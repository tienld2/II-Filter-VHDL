-------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   15:34:34 09/05/2013
-- Design Name:   
-- Module Name:   /home/nick/polyDecimDemodFilter2/polyDecimDemodFilter2_Top_tb.vhd
-- Project Name:  polyDecimDemodFilter2
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: polyDecimDemodFilter2_Top
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
use IEEE.std_logic_misc.all;
use IEEE.std_logic_unsigned.all;
use IEEE.MATH_REAL.all;


ENTITY polyDecimDemodFilter2_Top_tb IS
END polyDecimDemodFilter2_Top_tb;
 
ARCHITECTURE behavior OF polyDecimDemodFilter2_Top_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT polyDecimDemodFilter2_Top
    PORT(
      clk : in std_logic;
      clk_enable : in std_logic;
      max_count : in unsigned(3 downto 0);
      rst : in std_logic;
      tValidIn_Array : in std_logic_vector(15 downto 0) ;
      runSignals : in std_logic_vector(15 downto 0);
      reloadFIRCoefData : std_logic_vector(15 downto 0) ;
      phaseInc : in std_logic_vector(15 downto 0);
      accCoefs : in std_logic_vector(31 downto 0) ;
      trigger_array     : in std_logic_vector(4 downto 0) ;
      -- -------------------------------------------------
      -- temporary signals -------------------------------
      datatoDemodTop    : out std_logic_vector(19 downto 0) ;
      dataOutFromDemodRe  : out std_logic_vector(35 downto 0) ;
      dataOutFromDemodIm  : out std_logic_vector(35 downto 0) ;
      mulOutput       : out std_logic_vector(79 downto 0) ;
      blockRamOutput    : out std_logic_vector(31 downto 0) ;
      iirFilterTmp : out std_logic_vector(39 downto 0) ;
      -- temporary signals -------------------------------
      -- -------------------------------------------------
      inputSignal : in std_logic_vector(15 downto 0) ;
      outputDataRe : out std_logic_vector(19 downto 0) ;
      outputDataIm : out std_logic_vector(19 downto 0) ;
      acc : out std_logic_vector(99 downto 0)         );
    END COMPONENT;


   --Inputs
   signal clk : std_logic := '0';
   signal clk_enable : std_logic := '0';
   signal clk_div : std_logic := '0';                         --   (samplingFreq / decimFactor) / 2
   signal max_count : unsigned(3 downto 0) := b"0001";        --   (100 MHz      / 4          ) / 2 = 12500000 
   signal rst : std_logic := '0';
   signal tValidIn_Array : std_logic_vector(15 downto 0) := (others => '0');
   signal runSignals : std_logic_vector(15 downto 0) := (others => '0');
   signal reloadFIRCoefData : std_logic_vector(15 downto 0) := (others => '0');
   signal phaseInc : std_logic_vector(15 downto 0) := (others => '0');
   signal inputSignal : std_logic_vector(15 downto 0) := (others => '0');
   signal accCoefs : std_logic_vector(31 downto 0) ;
   signal trigger_array : std_logic_vector(4 downto 0) ;
   -- -------------------------------------------------
   -- temporary signals -------------------------------
   signal datatoDemodTop : std_logic_vector(19 downto 0) := (others => '0');
   signal dataOutFromDemodRe : std_logic_vector(35 downto 0) := (others => '0');
   signal dataOutFromDemodIm  : std_logic_vector(35 downto 0) := (others => '0');
   signal mulOutput : std_logic_vector(79 downto 0) ;
   signal blockRamOutput : std_logic_vector(31 downto 0) ;
   signal iirFilterTmp : std_logic_vector(39 downto 0) ;
   -- temporary signals -------------------------------
   -- -------------------------------------------------


  -- Constants
  constant inputSize : integer := 4001;
  constant coefSize : integer := 4095;

	--Outputs
 signal outputDataRe : std_logic_vector(19 downto 0);
 signal outputDataIm : std_logic_vector(19 downto 0);
 signal acc : std_logic_vector(99 downto 0) ;

 -- Clock period definitions
 constant clk_period : time := 10 ns;
 constant clk_enable_period : time := 10 ns;

  -- clock divided clock:
  signal clk_div_counter : integer := 0;
  signal clk_div_temp : std_logic := '1';

  -- padding for outputs
  signal padding : std_logic_vector(13 downto 0) := (others => '0');
  signal accReLSB, accImLSB : std_logic_vector(31 downto 0) ;


  type input_array is array (0 to inputSize) of std_logic_vector(15 downto 0) ;
  type input_array32 is array (inputSize downto 0) of std_logic_vector(31 downto 0) ;
signal myCosine : input_array :=(x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000");
     -- signal myCoef : input_array32 :=(x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");
signal myCoef : input_array32 := (others => x"00007fff");

BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: polyDecimDemodFilter2_Top PORT MAP (
          clk => clk,
          clk_enable => clk_enable,
          max_count => max_count,
          rst => rst,
          tValidIn_Array => tValidIn_Array,
          runSignals => runSignals,
          reloadFIRCoefData => reloadFIRCoefData,
          phaseInc => phaseInc,
          inputSignal => inputSignal,
          accCoefs => accCoefs,
          trigger_array => trigger_array,
          -- -------------------------------------------------
          -- temporary signals -------------------------------
          datatoDemodTop => datatoDemodTop,
          dataOutFromDemodRe => dataOutFromDemodRe,
          dataOutFromDemodIm => dataOutFromDemodIm,
          mulOutput => mulOutput,
          blockRamOutput => blockRamOutput,
          iirFilterTmp => iirFilterTmp,
          -- temporary signals -------------------------------
          -- -------------------------------------------------
          outputDataRe => outputDataRe,
          outputDataIm => outputDataIm,
          acc => acc
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 
   clk_enable_process :process
   begin
		clk_enable <= '0';
		wait for clk_enable_period/2;
		clk_enable <= '1';
		wait for clk_enable_period/2;
   end process;


   -- ------------------------------------------------------------------------------------------------------
   --                                       temporary signals 
   -- ------------------------------------------------------------------------------------------------------
   output_filedatatoDemodTop : entity work.file_writer 
   generic map( 
     dataWidth => 20,
     wordWidth => 1,
     -- dataFrac => 15,
     fileName => "/home/nick/polyDecimDemodFilter2/dataFromFIRFilteroutput10MHz.dat"
   )
   port map( 
     reset => rst,
     clk => clk_div,
     enable => tValidIn_Array(0),
     data => datatoDemodTop,
     data_valid => tValidIn_Array(0)
   );

   output_filedataDemodReoutput : entity work.file_writer 
   generic map( 
     dataWidth => 20,
     wordWidth => 1,
     -- dataFrac => 15,
     fileName => "/home/nick/polyDecimDemodFilter2/dataDemodReoutput10MHz.dat"
   )
   port map( 
     reset => rst,
     clk => clk_div,
     enable => tValidIn_Array(0),
     data => dataOutFromDemodRe(30 downto 11),
     data_valid => tValidIn_Array(0)
   );

   output_filedataDemodImoutput : entity work.file_writer 
   generic map( 
     dataWidth => 20,
     wordWidth => 1,
     -- dataFrac => 15,
     fileName => "/home/nick/polyDecimDemodFilter2/dataDemodImoutput10MHz.dat"
   )
   port map( 
     reset => rst,
     clk => clk_div,
     enable => tValidIn_Array(0),
     data => dataOutFromDemodIm(30 downto 11),
     data_valid => tValidIn_Array(0)
   );
   -- ------------------------------------------------------------------------------------------------------
   -- ------------------------------------------------------------------------------------------------------



   -- clk for file writer from iir filters:
   my_clk_div : entity work.clk_div_top
    port map(
      max_count => max_count,
      clk_in => clk,
      rst => rst,
      clk_out => clk_div
    ) ;

  output_fileCos : entity work.file_writer 
  generic map( 
    dataWidth => 16,
    wordWidth => 1,
    -- dataFrac => 15,
    fileName => "/home/nick/polyDecimDemodFilter2/cosoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk,
    enable => tValidIn_Array(0),
    data => inputSignal,
    data_valid => tValidIn_Array(0)
  );



  output_fileiirreal : entity work.file_writer 
  generic map( 
    dataWidth => 20,
    wordWidth => 1,
    -- dataFrac => 15,
    fileName => "/home/nick/polyDecimDemodFilter2/dataIIRFilterReoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk_div,
    enable => tValidIn_Array(0),
    data => iirFilterTmp(19 downto 0),
    data_valid => tValidIn_Array(0)
  );


  output_fileiirimag : entity work.file_writer 
  generic map( 
    dataWidth => 20,
    wordWidth => 1,
    -- dataFrac => 15,
    fileName => "/home/nick/polyDecimDemodFilter2/dataIIRFilterImoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk_div,
    enable => tValidIn_Array(0),
    data => iirFilterTmp(39 downto 20),
    data_valid => tValidIn_Array(0)
  );

  -- ------------------------------------------------------------------------------------------------------
  --                        plotted with plotChannelizer.py
  -- ------------------------------------------------------------------------------------------------------

  -- output_fileRe : entity work.file_writer 
  -- generic map( 
  --   dataWidth => 20,
  --   wordWidth => 1,
  --   -- dataFrac => 10,
  --   fileName => "/home/nick/polyDecimDemodFilter2/polyDecimDemodFilter2Reoutput10MHz.dat"
  -- )
  -- port map( 
  --   reset => rst,
  --   clk => clk_div,
  --   enable => '1',
  --   data => outputDataRe,
  --   data_valid => '1'
  -- );

  -- output_fileIm : entity work.file_writer 
  -- generic map( 
  --   dataWidth => 20,
  --   wordWidth => 1,
  --   -- dataFrac => 10,
  --   fileName => "/home/nick/polyDecimDemodFilter2/polyDecimDemodFilter2Imoutput10MHz.dat"
  -- )
  -- port map( 
  --   reset => rst,
  --   clk => clk_div,
  --   enable => '1',
  --   data => outputDataIm,
  --   data_valid => '1'
  -- );

  -- ------------------------------------------------------------------------------------------------------
  -- ------------------------------------------------------------------------------------------------------

accReLSB <= padding & acc(17 downto 0);
accImLSB <= padding & acc(67 downto 50);


-- Bottom 32 bits of output
output_filemacReLSB : entity work.file_writer 
generic map( 
  dataWidth => 32,
  wordWidth => 1,
  -- dataFrac => 10,
  fileName => "/home/nick/polyDecimDemodFilter2/polyDecimDemodFilter2ReLSBoutput10MHz.dat"
)
port map( 
  reset => rst,
  clk => clk_div,
  enable => trigger_array(2),
  data => acc(31 downto 0),
  data_valid => trigger_array(2)
);

output_filemacImLSB : entity work.file_writer 
  generic map( 
    dataWidth => 32,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/polyDecimDemodFilter2/polyDecimDemodFilter2ImLSBoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk_div,
    enable => trigger_array(2),
    data => acc(81 downto 50),
    data_valid => trigger_array(2)
  );

-- Top 18 bits of output
output_filemacReMSB : entity work.file_writer 
  generic map( 
    dataWidth => 18,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/polyDecimDemodFilter2/polyDecimDemodFilter2ReMSBoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk_div,
    enable => trigger_array(2),
    data => acc(49 downto 32),
    data_valid => trigger_array(2)
  );

output_filemacImMSB : entity work.file_writer 
  generic map( 
    dataWidth => 18,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/polyDecimDemodFilter2/polyDecimDemodFilter2ImMSBoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk_div,
    enable => trigger_array(2),
    data => acc(99 downto 82),
    data_valid => trigger_array(2)
  );


  output_fileWindow : entity work.file_writer 
  generic map( 
    dataWidth => 32,
    wordWidth => 1,
    -- dataFrac => 15,
    fileName => "/home/nick/polyDecimDemodFilter2/dataMULwindowoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk_div,
    enable => trigger_array(2),
    data => blockRamOutput,
    data_valid => trigger_array(2)
  );

  -- temporary signals ---------------------------------------------------
output_filemulRe : entity work.file_writer 
  generic map( 
    dataWidth => 36,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/polyDecimDemodFilter2/dataMULReoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk_div,
    enable => trigger_array(2),
    data => mulOutput(35 downto 0),
    data_valid => trigger_array(2)
  );

output_filemulIm : entity work.file_writer 
  generic map( 
    dataWidth => 36,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/polyDecimDemodFilter2/dataMULImoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk_div,
    enable => trigger_array(2),
    data => mulOutput(75 downto 40),
    data_valid => trigger_array(2)
  );
-- temporary signals ---------------------------------------------------





   -- Stimulus process
   stim_proc: process
   begin		

      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;

      -- Initialize all inputs, then reset
      -- acc <= (others => '0');
      trigger_array <= (others => '0');
      runSignals <= (others => '0');
      accCoefs <= (others => '0');

      -- insert, stimulus here 
      -- pulse the reset line:
      rst <= '1'; wait until (rising_edge(clk));
      wait for clk_period*20;
      rst <= '0'; wait until (rising_edge(clk));
      report "System reset with global signal rst.\n";

      report "Coefficients initialized to 0...\n";
      -- mac block ram instructions 
      -- -----------------------------------------------------------
      -- load coefficient block ram:
      trigger_array(1) <= '1'; wait until (rising_edge(clk)); 
      report "Setting write_en to populate block ram with coefs...";
      for i in 0 to inputSize loop
        accCoefs <= myCoef(i); wait until (rising_edge(clk)); 
      end loop;
      report "Coefficients loaded into block ram.";
      trigger_array(1) <= '0'; wait until (rising_edge(clk)); 

      -- feed data into polyDecimator, start filtering:
      tValidIn_Array(0) <= '1'; wait until (rising_edge(clk));
      runSignals(0) <= '1'; wait until (rising_edge(clk));
      report "polyDecimator triggered, transmitting data to filter now...\n";

      tValidIn_Array(1) <= '1';
      trigger_array(2) <= '1'; 
            phaseInc <= x"147A"; wait until (rising_edge(clk));           
            -- phaseInc <= x"0000"; wait until (rising_edge(clk));           
      report "Setting phaseInc to x'147A', initiating demodulator...\n";

      for i in 0 to inputSize loop
        inputSignal <= myCosine(i); wait until (rising_edge(clk)); 
      end loop;


      -- start reading input data and start accumulating:
      report "\nStarting multiply-accumulator...";
 
      report "Finished reading input data.";

      runSignals <= (others => '0');
      report "Finished processing.";

      wait;
   end process;

END;
