--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   09:45:26 09/23/2013
-- Design Name:   
-- Module Name:   /home/nick/mac16/mac16_top_tb.vhd
-- Project Name:  mac16
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: mac16_top
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.ALL;
use IEEE.std_logic_misc.all;
use IEEE.std_logic_unsigned.all;

 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY mac16_top_tb IS
END mac16_top_tb;
 
ARCHITECTURE behavior OF mac16_top_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT mac16_top
    PORT(
      clk_in        : in std_logic;
      clk         : in std_logic;
      clk_en        : in std_logic;
      rst         : in std_logic;
      trigger_array     : in std_logic_vector(4 downto 0) ;
      coefDataIn      : in std_logic_vector(31 downto 0) ;
      iirData       : in std_logic_vector(39 downto 0) ;
      -- tempory signals --------------------------------------
      mulOutput       : out std_logic_vector(79 downto 0) ;
      blockRamOutput  : out std_logic_vector(31 downto 0) ;
      -- tempory signals --------------------------------------
      acc         : out std_logic_vector(95 downto 0)         );
    END COMPONENT;
    

   --Inputs
   signal clk_in : std_logic := '0';
   signal clk : std_logic := '0';
   signal clk_en : std_logic := '0';
   signal rst : std_logic := '0';
   signal trigger_array : std_logic_vector(4 downto 0) := (others => '0');
   signal coefDataIn : std_logic_vector(31 downto 0) := (others => '0');
   signal iirData : std_logic_vector(39 downto 0) := (others => '0');

   

 	--Outputs
   signal acc : std_logic_vector(95 downto 0);
  
  -- tempory signals --------------------------------------
  signal mulOutput : std_logic_vector(79 downto 0) ;
  signal blockRamOutput  : std_logic_vector(31 downto 0) ;
  -- tempory signals --------------------------------------
  

   -- Clock period definitions
   constant clk_in_period : time := 40 ns;
   constant clk_period : time := 10 ns;
   constant clk_en_period : time := 10 ns;

   constant inputSize : integer := 4095;

   type input_array40 is array (inputSize downto 0) of std_logic_vector(39 downto 0) ;
   type input_array32 is array (inputSize downto 0) of std_logic_vector(31 downto 0) ;
   signal myCosine : input_array40 :=(x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"00FFFE803F",x"00FFFF7F68",x"0000008098",x"0000017FC1",x"00000278DD",x"00000367FE",x"000004495F",x"0000051971",x"000005D4EC",x"00000678DD",x"00000702AC",x"000007702D",x"000007BFA7",x"000007EFD8",x"000007FFFF",x"000007EFD8",x"000007BFA7",x"000007702D",x"00000702AC",x"00000678DD",x"000005D4EC",x"0000051971",x"000004495F",x"00000367FE",x"00000278DD",x"0000017FC1",x"0000008098",x"00FFFF7F68",x"00FFFE803F",x"00FFFD8723",x"00FFFC9802",x"00FFFBB6A1",x"00FFFAE68F",x"00FFFA2B14",x"00FFF98723",x"00FFF8FD54",x"00FFF88FD3",x"00FFF84059",x"00FFF81028",x"00FFF80001",x"00FFF81028",x"00FFF84059",x"00FFF88FD3",x"00FFF8FD54",x"00FFF98723",x"00FFFA2B14",x"00FFFAE68F",x"00FFFBB6A1",x"00FFFC9802",x"00FFFD8723",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"00FFF82448",x"00FFF8040C",x"00FFF8040C",x"00FFF82448",x"00FFF8643E",x"00FFF8C2EB",x"00FFF93ED2",x"00FFF9D5FE",x"00FFFA860D",x"00FFFB4C38",x"00FFFC255F",x"00FFFD0E16",x"00FFFE02B0",x"00FFFEFF52",x"0000000000",x"00000100AE",x"000001FD50",x"000002F1EA",x"000003DAA1",x"000004B3C8",x"00000579F3",x"0000062A02",x"000006C12E",x"0000073D15",x"0000079BC2",x"000007DBB8",x"000007FBF4",x"000007FBF4",x"000007DBB8",x"0000079BC2",x"0000073D15",x"000006C12E",x"0000062A02",x"00000579F3",x"000004B3C8",x"000003DAA1",x"000002F1EA",x"000001FD50",x"00000100AE",x"0000000000",x"00FFFEFF52",x"00FFFE02B0",x"00FFFD0E16",x"00FFFC255F",x"00FFFB4C38",x"00FFFA860D",x"00FFF9D5FE",x"00FFF93ED2",x"00FFF8C2EB",x"00FFF8643E",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000",x"0000000000");
   signal myCoef : input_array32 :=(x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

 
BEGIN
 
  
	-- Instantiate the Unit Under Test (UUT)
   uut: mac16_top PORT MAP (
          clk_in => clk_in,
          clk => clk,
          clk_en => clk_en,
          rst => rst,
          trigger_array => trigger_array,
          coefDataIn => coefDataIn,
          iirData => iirData,
          -- tempory signals --------------------------------------
          mulOutput => mulOutput,
          blockRamOutput => blockRamOutput,
          -- tempory signals --------------------------------------
          acc => acc
        );

   -- Clock process definitions
   clk_in_process :process
   begin
		clk_in <= '0';
		wait for clk_in_period/2;
		clk_in <= '1';
		wait for clk_in_period/2;
   end process;
 
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 
   clk_en_process :process
   begin
		clk_en <= '0';
		wait for clk_en_period/2;
		clk_en <= '1';
		wait for clk_en_period/2;
   end process;
 
  output_fileCosRe : entity work.file_writer 
  generic map( 
    dataWidth => 20,
    wordWidth => 1,
    -- dataFrac => 15,
    fileName => "/home/nick/mac16/cosoutputRe10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk,
    enable => trigger_array(1),
    data => iirData(19 downto 0),
    data_valid => trigger_array(1)
  );

  output_fileCosIm : entity work.file_writer 
  generic map( 
    dataWidth => 20,
    wordWidth => 1,
    -- dataFrac => 15,
    fileName => "/home/nick/mac16/cosoutputIm10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk,
    enable => trigger_array(1),
    data => iirData(39 downto 20),
    data_valid => trigger_array(1)
  );

  output_fileWindow : entity work.file_writer 
  generic map( 
    dataWidth => 32,
    wordWidth => 1,
    -- dataFrac => 15,
    fileName => "/home/nick/mac16/dataMULwindowoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk,
    enable => trigger_array(2),
    data => blockRamOutput,
    data_valid => trigger_array(2)
  );


-- temporary signals ---------------------------------------------------
output_filemulRe : entity work.file_writer 
  generic map( 
    dataWidth => 36,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/mac16/dataMULReoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk,
    enable => trigger_array(2),
    data => mulOutput(35 downto 0),
    data_valid => trigger_array(2)
  );

output_filemulIm : entity work.file_writer 
  generic map( 
    dataWidth => 36,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/mac16/dataMULImoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk,
    enable => trigger_array(2),
    data => mulOutput(75 downto 40),
    data_valid => trigger_array(2)
  );
-- temporary signals ---------------------------------------------------

  output_filemacRe : entity work.file_writer 
  generic map( 
    dataWidth => 48,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/mac16/mac16Reoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk,
    enable => trigger_array(2),
    data => acc(47 downto 0),
    data_valid => trigger_array(2)
  );

output_filemacIm : entity work.file_writer 
  generic map( 
    dataWidth => 48,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/mac16/mac16Imoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk,
    enable => trigger_array(2),
    data => acc(95 downto 48),
    data_valid => trigger_array(2)
  );



   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_in_period*10;

      -- insert stimulus here 
      
      -- pump rst lines:
      rst <= '1'; wait until (rising_edge(clk));
      wait for clk_period*4;
      rst <= '0'; wait until (rising_edge(clk));
      report "System reset with global signal rst.\n";

      -- trigger block ram coef writing:
      trigger_array(1) <= '1'; wait until (rising_edge(clk)); 
      report "Setting write_en to populate block ram with coefs...";
      for i in 0 to inputSize loop
        coefDataIn <= myCoef(i); wait until (rising_edge(clk)); 
      end loop;
      report "Coefficients loaded into block ram.";
      

      -- start reading input data and start accumulating:
      trigger_array(2) <= '1'; 
      report "\nStarting multiply-accumulator...";
      for i in 0 to inputSize loop
        iirData <= myCosine(i); wait until (rising_edge(clk)); 
      end loop;
      report "Finished reading input data.";

      trigger_array <= (others => '0'); 
      report "\nFinished Processing.";


      wait;
   end process;

END;
