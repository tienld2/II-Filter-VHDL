-- Copyright 2010 by Innovative Integration Inc., All Rights Reserved.
--******************************************************************************
--* Design Name: ii_dac_bitslip
--*
--* @li Target Device: any
--* @li Tool versions: ISE 12.3
--*
--*     @short DAC output alignment control with external sync
--*
--* Description:
--*
--*   This module adjusts the DAC data latency based on the ext_sync_phase
--*   value latched when an ext_sync occurs to maintain a fixed delay between
--*   the ext_sync and the DAC output.
--*
--*
--*   @port dac_clk_bufr    : input, regional clock generated by dividing
--*                                  dac_clk_in using BUFR
--*   @port trig_clk_phase  : input, latched clock phase on trigger
--*   @port dac_dual_ch     : input, DAC is in dual channel mode
--*   @port dac_dll_bypass  : input, DAC dll is bypassed
--*   @port dac_shift_cnt   : input, DAC output shift count
--*   @port ext_sync_phase  : input, external sync phase
--*   @port raw_sync        : input, raw DAC sync
--*   @port raw_data        : input, raw DAC data
--*   @port algnd_sync      :output, aligned DAC sync
--*   @port algnd_data      :output, aligned DAC data
--*
--*      @author Innovative Integration
--*      @version 1.0
--*      @date Created 11/23/10
--*
--******************************************************************************
--/

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ii_dac_bitslip is
  port (
    -- clock
    dac_clk_bufr         : in  std_logic;

    -- control
    trig_clk_phase       : in  std_logic;
    dac_dual_ch          : in  std_logic;
    dac_dll_bypass       : in  std_logic;
    dac_shift_cnt        : in  std_logic_vector(3 downto 0);
    ext_sync_phase       : in  std_logic_vector(1 downto 0);

    -- raw DAC data
    raw_sync             : in  std_logic;
    raw_data             : in  std_logic_vector(63 downto 0);

    -- aligned DAC data
    algnd_sync           : out std_logic_vector(3 downto 0);
    algnd_data           : out std_logic_vector(63 downto 0)
  );
end ii_dac_bitslip;

architecture arch of ii_dac_bitslip is

  signal es_shift_cnt         : unsigned(2 downto 0);
  signal trig_lat             : integer;
  signal bitslip_cnt          : unsigned(4 downto 0);
  signal raw_sync_1d          : std_logic;
  signal raw_sync_2d          : std_logic;
  signal raw_sync_3d          : std_logic;
  signal raw_sync_4d          : std_logic;
  signal raw_sync_5d          : std_logic;
  signal raw_sync_6d          : std_logic;
  signal raw_data_1d          : std_logic_vector(63 downto 0);
  signal raw_data_2d          : std_logic_vector(63 downto 0);
  signal raw_data_3d          : std_logic_vector(63 downto 0);
  signal raw_data_4d          : std_logic_vector(63 downto 0);
  signal raw_data_5d          : std_logic_vector(63 downto 0);
  signal raw_data_6d          : std_logic_vector(63 downto 0);

begin

  -- Calculate the shift amount for different configurations
  process (dac_clk_bufr)
  begin
    if (rising_edge(dac_clk_bufr)) then
      if (dac_dual_ch = '0' and dac_dll_bypass = '0') then
        es_shift_cnt <= '0' & unsigned(ext_sync_phase);
      elsif (dac_dual_ch = '1' and dac_dll_bypass = '1') then
        case (ext_sync_phase) is
          when "00" =>
            es_shift_cnt <= "000";
          when others =>
            es_shift_cnt <= "100";
        end case;
      else
        case (ext_sync_phase) is
          when "01" | "10"=>
            es_shift_cnt <= "010";
          when "11" =>
            es_shift_cnt <= "100";
          when others =>
            es_shift_cnt <= "000";
        end case;
      end if;
    end if;
  end process;

  -- Delay required when the DLL is disabled
  trig_lat <= 4 when (trig_clk_phase = '1' and dac_dll_bypass = '1') else
              0;

  -- Add up the three shift values to make up the final bitslip count
  process (dac_clk_bufr)
  begin
    if (rising_edge(dac_clk_bufr)) then
      bitslip_cnt <= to_unsigned(trig_lat,5) + resize(es_shift_cnt,5) +
                     resize(unsigned(dac_shift_cnt),5);
    end if;
  end process;

  -- Pipeline raw_sync and raw_data
  process (dac_clk_bufr)
  begin
    if (rising_edge(dac_clk_bufr)) then
      raw_sync_1d <= raw_sync;
      raw_sync_2d <= raw_sync_1d;
      raw_sync_3d <= raw_sync_2d;
      raw_sync_4d <= raw_sync_3d;
      raw_sync_5d <= raw_sync_4d;
      raw_sync_6d <= raw_sync_5d;
      raw_data_1d <= raw_data;
      raw_data_2d <= raw_data_1d;
      raw_data_3d <= raw_data_2d;
      raw_data_4d <= raw_data_3d;
      raw_data_5d <= raw_data_4d;
      raw_data_6d <= raw_data_5d;
    end if;
  end process;

  -- Delay logic
  process (dac_clk_bufr)
  begin
    if (rising_edge(dac_clk_bufr)) then
      case (bitslip_cnt) is
        when "00000" =>
          algnd_sync <= raw_sync_1d & raw_sync_1d & raw_sync_1d & raw_sync_1d;
          algnd_data <= raw_data_1d;
        when "00001" =>
          algnd_sync <= raw_sync_1d & raw_sync_1d & raw_sync_1d & raw_sync_2d;
          algnd_data <= raw_data_1d(47 downto 0) & raw_data_2d(63 downto 48);
        when "00010" =>
          algnd_sync <= raw_sync_1d & raw_sync_1d & raw_sync_2d & raw_sync_2d;
          algnd_data <= raw_data_1d(31 downto 0) & raw_data_2d(63 downto 32);
        when "00011" =>
          algnd_sync <= raw_sync_1d & raw_sync_2d & raw_sync_2d & raw_sync_2d;
          algnd_data <= raw_data_1d(15 downto 0) & raw_data_2d(63 downto 16);
        when "00100" =>
          algnd_sync <= raw_sync_2d & raw_sync_2d & raw_sync_2d & raw_sync_2d;
          algnd_data <= raw_data_2d;
        when "00101" =>
          algnd_sync <= raw_sync_2d & raw_sync_2d & raw_sync_2d & raw_sync_3d;
          algnd_data <= raw_data_2d(47 downto 0) & raw_data_3d(63 downto 48);
        when "00110" =>
          algnd_sync <= raw_sync_2d & raw_sync_2d & raw_sync_3d & raw_sync_3d;
          algnd_data <= raw_data_2d(31 downto 0) & raw_data_3d(63 downto 32);
        when "00111" =>
          algnd_sync <= raw_sync_2d & raw_sync_3d & raw_sync_3d & raw_sync_3d;
          algnd_data <= raw_data_2d(15 downto 0) & raw_data_3d(63 downto 16);
        when "01000" =>
          algnd_sync <= raw_sync_3d & raw_sync_3d & raw_sync_3d & raw_sync_3d;
          algnd_data <= raw_data_3d;
        when "01001" =>
          algnd_sync <= raw_sync_3d & raw_sync_3d & raw_sync_3d & raw_sync_4d;
          algnd_data <= raw_data_3d(47 downto 0) & raw_data_4d(63 downto 48);
        when "01010" =>
          algnd_sync <= raw_sync_3d & raw_sync_3d & raw_sync_4d & raw_sync_4d;
          algnd_data <= raw_data_3d(31 downto 0) & raw_data_4d(63 downto 32);
        when "01011" =>
          algnd_sync <= raw_sync_3d & raw_sync_4d & raw_sync_4d & raw_sync_4d;
          algnd_data <= raw_data_3d(15 downto 0) & raw_data_4d(63 downto 16);
        when "01100" =>
          algnd_sync <= raw_sync_4d & raw_sync_4d & raw_sync_4d & raw_sync_4d;
          algnd_data <= raw_data_4d;
        when "01101" =>
          algnd_sync <= raw_sync_4d & raw_sync_4d & raw_sync_4d & raw_sync_5d;
          algnd_data <= raw_data_2d(47 downto 0) & raw_data_3d(63 downto 48);
        when "01110" =>
          algnd_sync <= raw_sync_4d & raw_sync_4d & raw_sync_5d & raw_sync_5d;
          algnd_data <= raw_data_4d(31 downto 0) & raw_data_5d(63 downto 32);
        when "01111" =>
          algnd_sync <= raw_sync_4d & raw_sync_5d & raw_sync_5d & raw_sync_5d;
          algnd_data <= raw_data_4d(15 downto 0) & raw_data_5d(63 downto 16);
        when "10000" =>
          algnd_sync <= raw_sync_5d & raw_sync_5d & raw_sync_5d & raw_sync_5d;
          algnd_data <= raw_data_5d;
        when "10001" =>
          algnd_sync <= raw_sync_5d & raw_sync_5d & raw_sync_5d & raw_sync_6d;
          algnd_data <= raw_data_5d(47 downto 0) & raw_data_6d(63 downto 48);
        when "10010" =>
          algnd_sync <= raw_sync_5d & raw_sync_5d & raw_sync_6d & raw_sync_6d;
          algnd_data <= raw_data_5d(31 downto 0) & raw_data_6d(63 downto 32);
        when "10011" =>
          algnd_sync <= raw_sync_5d & raw_sync_6d & raw_sync_6d & raw_sync_6d;
          algnd_data <= raw_data_5d(15 downto 0) & raw_data_6d(63 downto 16);
        when "10100" =>
          algnd_sync <= raw_sync_6d & raw_sync_6d & raw_sync_6d & raw_sync_6d;
          algnd_data <= raw_data_6d;
        when others =>
      end case;
    end if;
  end process;

end arch;
