-- Copyright 2010 by Innovative Integration Inc., All Rights Reserved.
--******************************************************************************
--* Design Name: ii_dac5682z_intf
--*
--* @li Target Device: Virtex-6
--* @li Tool versions: ISE 13.2
--*
--*     @short D/A interface for TI DAC5682Z
--*
--* Description:
--*
--*   This file is the interface to DAC5682z. It receives streaming data
--*   or test data (if test enabled) over a 64 bit parallel bus at sys_clk
--*   domain and stores them in a FIFO.
--*   When triggered, the FIFO is read and the read data is routed to the
--*   DAC physical layer interface that serializes the slow rate parallel
--*   input into a serial stream at a higher rate at the DAC interface.
--*
--*
--*   @port srst            : input, synchronous active high reset
--*   @port dac_reset       : input, synchronous active high DAC reset
--*                                  @sys_clk domain
--*   @port sys_clk         : input, system clock
--*   @port dac_clk_bufio   :output, IO clock
--*   @port dac_clk_bufr    :output, regional clock generated by dividing
--*                                  dac_clk_in using BUFR
--*   @port dac_run         : input, enable DAC
--*   @port test_en         : input, test enable
--*   @port test_mode       : input, test mode select
--*   @port phase_inc_wr    : input, phase increment write strobe
--*   @port phase_inc       : input, phase increment
--*   @port dac_dual_ch     : input, DAC is in dual channel mode
--*   @port dac_dll_bypass  : input, DAC dll is bypassed
--*   @port dac_a_gain      : input, DAC-A gain correction coefficient (2's complement)
--*   @port dac_a_offset    : input, DAC-A offset correction coefficient (2's complement)
--*   @port dac_b_gain      : input, DAC-B gain correction coefficient (2's complement)
--*   @port dac_b_offset    : input, DAC-B offset correction coefficient (2's complement)
--*   @port ext_sync        : input, external sync (trigger) input
--*   @port ext_sync_phase  : input, external sync phase
--*   @port sw_trig         : input, software trigger input
--*   @port window_size     : input, number of points in a frame count
--*   @port trigger_mode    : input, trigger mode
--*   @port dac_trigger_en  :output, DAC trigger window is enabled
--*   @port dac_trig_alrt   :output, DAC trigger occurred
--*   @port underflow       :output, fifo underflow occurred
--*   @port din_wr          : input, data write strobe
--*   @port din             : input, data input
--*   @port fifo_rdy        :output, DAC fifo ready (with room)
--*   @port idelayctrl_rst  : input, synchronous active high reset, must
--*                                  be set for at least 50ns after configuration
--*                                  and ref_clk200 stabilized
--*   @port ref_clk200      : input, reference clock 200MHz needed by IDELAYCTRL
--*   @port dac_cal_en      : input, enable latency calibration
--*   @port dac_cal0_done   :output, DAC calibration 0 done
--*   @port dac_cal1_done   :output, DAC calibration 1 done
--*   @port dac_iodly_cnt   :output, DAC iodelay tap count
--*   @port dac_shift_cnt   :output, DAC output shift count
--*   @port dac_dig_p       : input, DAC digitized output differential pair (side-P)
--*   @port dac_dig_n       : input, DAC digitized output differential pair (side-N)
--*   @port dac_clk_in_p    : input, DAC clock differential pair (side-P)
--*   @port dac_clk_in_n    : input, DAC clock differential pair (side-N)
--*   @port dac_clk_out_p   :output, forwarded DAC clock differential pair (side-P)
--*   @port dac_clk_out_n   :output, forwarded DAC clock differential pair (side-N)
--*   @port sync_out_p      :output, DAC SYNC differential pair (side-P)
--*   @port sync_out_n      :output, DAC SYNC differential pair (side-N)
--*   @port sync2_out_p     :output, a copy of DAC SYNC differential pair (side-P)
--*   @port sync2_out_n     :output, a copy of DAC SYNC differential pair (side-N)
--*   @port data_out_p      :output, DAC Data differential pair (side-P) (16 bits)
--*   @port data_out_n      :output, DAC Data differential pair (side-N) (16 bits)
--*
--*      @author Innovative Integration
--*      @version 1.0
--*      @date Created 11/23/10
--*
--******************************************************************************
--/

library ieee;
use ieee.std_logic_1164.all;

entity ii_dac5682z_intf is
  port (
    -- Resets and clocks
    srst                 : in  std_logic;
    dac_reset            : in  std_logic;
    sys_clk              : in  std_logic;
    dac_clk_bufio        : out std_logic;
    dac_clk_bufr         : out std_logic;

    -- Control
    dac_run              : in  std_logic;
    test_en              : in  std_logic;
    test_mode            : in  std_logic_vector(2 downto 0);
    phase_inc_wr         : in  std_logic;
    phase_inc            : in  std_logic_vector(31 downto 0);
    dac_dual_ch          : in  std_logic;
    dac_dll_bypass       : in  std_logic;
    dac_a_gain           : in  std_logic_vector(17 downto 0);
    dac_a_offset         : in  std_logic_vector(15 downto 0);
    dac_b_gain           : in  std_logic_vector(17 downto 0);
    dac_b_offset         : in  std_logic_vector(15 downto 0);

    -- External Sync and trigger interface
    ext_sync             : in  std_logic;
    ext_sync_phase       : in  std_logic_vector(1 downto 0);
    sw_trig              : in  std_logic;
    window_size          : in  std_logic_vector(23 downto 0);
    trigger_mode         : in  std_logic_vector(2 downto 0);
    dac_trigger_en       : out std_logic;

    -- Alerts
    dac_trig_alrt        : out std_logic;
    underflow            : out std_logic;

    -- Data fifo interface
    din_wr               : in  std_logic;
    din                  : in  std_logic_vector(63 downto 0);
    fifo_rdy             : out std_logic;

    -- reference clock
    idelayctrl_rst       : in  std_logic;
    ref_clk200           : in  std_logic;

    -- Latency calibration control and status
    dac_cal_en           : in  std_logic;
    dac_cal0_done        : out std_logic;
    dac_cal1_done        : out std_logic;
    dac_iodly_cnt        : out std_logic_vector(4 downto 0);
    dac_shift_cnt        : out std_logic_vector(3 downto 0);

    -- DAC output digitizer interface
    dac_dig_p            : in  std_logic;
    dac_dig_n            : in  std_logic;

    -- DAC interface signals
    dac_clk_in_p         : in  std_logic;
    dac_clk_in_n         : in  std_logic;
    dac_clk_out_p        : out std_logic;
    dac_clk_out_n        : out std_logic;
    sync_out_p           : out std_logic;
    sync_out_n           : out std_logic;
    sync2_out_p          : out std_logic;
    sync2_out_n          : out std_logic;
    data_out_p           : out std_logic_vector(15 downto 0);
    data_out_n           : out std_logic_vector(15 downto 0)
  );
end ii_dac5682z_intf;

architecture arch of ii_dac5682z_intf is

  component ii_offgain
    port (
      srst                 : in  std_logic;
      clk                  : in  std_logic;
      gain                 : in  std_logic_vector(17 downto 0);
      offset               : in  std_logic_vector(15 downto 0);
      ce                   : in  std_logic;
      din                  : in  std_logic_vector(15 downto 0);
      data_vld             : out std_logic;
      dout                 : out std_logic_vector(15 downto 0)
    );
  end component;

  component ii_trigger
    generic (
      SAMPLES_PER_CLK      : integer := 1
    );
    port (
      reset                : in  std_logic;
      clk                  : in  std_logic;
      ce                   : in  std_logic;
      ext_sync             : in  std_logic;
      sw_trig              : in  std_logic;
      trig_mode            : in  std_logic_vector(2 downto 0);
      frame_size           : in  std_logic_vector(23 downto 0);
      decimation_coeff     : in  std_logic_vector(11 downto 0);
      decimation_en        : out std_logic;
      trigger              : out std_logic;
      trigger_en           : out std_logic
    );
  end component;

  component ii_dac_bitslip
    port (
      -- clock
      dac_clk_bufr         : in  std_logic;

      -- control
      trig_clk_phase       : in  std_logic;
      dac_dual_ch          : in  std_logic;
      dac_dll_bypass       : in  std_logic;
      dac_shift_cnt        : in  std_logic_vector(3 downto 0);
      ext_sync_phase       : in  std_logic_vector(1 downto 0);

      -- raw DAC data
      raw_sync             : in  std_logic;
      raw_data             : in  std_logic_vector(63 downto 0);

      -- aligned DAC data
      algnd_sync           : out std_logic_vector(3 downto 0);
      algnd_data           : out std_logic_vector(63 downto 0)
    );
  end component;

  component ii_dac5682z_phy
    port (
      phy_rst              : in  std_logic;
      idelayctrl_rst       : in  std_logic;
      ref_clk200           : in  std_logic;
      dac_clk_bufio        : out std_logic;
      dac_clk_bufr         : out std_logic;
      dac_dll_bypass       : in  std_logic;

      -- Parallel data and output enable
      sync_in              : in  std_logic_vector(3 downto 0);
      data_in              : in  std_logic_vector(63 downto 0);

      -- DAC interface signals
      dac_clk_in_p         : in  std_logic;
      dac_clk_in_n         : in  std_logic;
      dac_clk_out_p        : out std_logic;
      dac_clk_out_n        : out std_logic;
      sync_out_p           : out std_logic;
      sync_out_n           : out std_logic;
      sync2_out_p          : out std_logic;
      sync2_out_n          : out std_logic;
      data_out_p           : out std_logic_vector(15 downto 0);
      data_out_n           : out std_logic_vector(15 downto 0)
    );
  end component;

  component ii_dac_lat_cal
    port (
      -- Reset and clocks
      dac_reset            : in  std_logic;
      fs_clk               : in  std_logic;
      fs_clkdiv2           : in  std_logic;

      -- Controls
      dac_cal_en           : in  std_logic;
      dac_run              : in  std_logic;
      dac_dual_ch          : in  std_logic;
      dac_dll_bypass       : in  std_logic;

      -- DAC output digitizer interface
      dac_dig_p            : in  std_logic;
      dac_dig_n            : in  std_logic;

      -- Outputs
      cal_trigger          : out std_logic;
      dac_cal0_done        : out std_logic;
      dac_cal1_done        : out std_logic;
      dac_iodly_cnt        : out std_logic_vector(4 downto 0);
      dac_shift_cnt        : out std_logic_vector(3 downto 0)
    );
  end component;

  component ii_dac_test_gen
    port (
      -- Reset and clock
      srst                 : in  std_logic;
      sys_clk              : in  std_logic;

      -- Control
      test_en              : in  std_logic;
      test_mode            : in  std_logic_vector(2 downto 0);
      phase_inc_wr         : in  std_logic;
      phase_inc            : in  std_logic_vector(31 downto 0);

      -- Data
      test_data_req        : in  std_logic;
      dout                 : out std_logic_vector(63 downto 0);
      valid                : out std_logic;
      pattern_test         : out std_logic
    );
  end component;

  component afifo_512x64_bram
    port (
      rst                  : in  std_logic;
      wr_clk               : in  std_logic;
      rd_clk               : in  std_logic;
      din                  : in  std_logic_vector(63 downto 0);
      wr_en                : in  std_logic;
      rd_en                : in  std_logic;
      dout                 : out std_logic_vector(63 downto 0);
      full                 : out std_logic;
      empty                : out std_logic;
      valid                : out std_logic;
      underflow            : out std_logic;
      prog_full            : out std_logic
    );
  end component;

  signal dac_rst_sreg         : std_logic_vector(3 downto 0);
  signal phy_rst              : std_logic;
  signal fifo_rst             : std_logic;
  signal selected_wr          : std_logic;
  signal selected_din         : std_logic_vector(63 downto 0);
  signal offgain_vld          : std_logic;
  signal offgain_dout         : std_logic_vector(63 downto 0);
  signal fifo_afull           : std_logic;
  signal fifo_afull_d         : std_logic;
  signal fifo_rdy_l           : std_logic;
  signal fifo_dout            : std_logic_vector(63 downto 0);
  signal fifo_dout_d          : std_logic_vector(63 downto 0);
  signal raw_data             : std_logic_vector(63 downto 0);
  signal fifo_underflow       : std_logic;
  signal fifo_underflow_d     : std_logic;
  signal fifo_underflow_dd    : std_logic;
  signal underflow_latch      : std_logic;
  signal underflow_latch_xdom : std_logic;
  signal underflow_latch_demet: std_logic;
  signal trigger              : std_logic;
  signal dac_clk_bufio_l      : std_logic;
  signal dac_clk_bufr_l       : std_logic;
  signal ph_en                : std_logic := '0';
  signal fifo_rden            : std_logic;
  signal fifo_dout_vld        : std_logic;
  signal fifo_dout_vld_d      : std_logic;
  signal fifo_dout_vld_dd     : std_logic;
  signal raw_sync             : std_logic;
  signal trigger_d            : std_logic;
  signal trigger_re           : std_logic;
  signal trigger_latch        : std_logic;
  signal trigger_latch_xdom   : std_logic;
  signal trigger_latch_demet  : std_logic;
  signal trig_clk_phase       : std_logic;
  signal offgain_0_2_gain     : std_logic_vector(17 downto 0);
  signal offgain_0_2_offset   : std_logic_vector(15 downto 0);
  signal offgain_1_3_gain     : std_logic_vector(17 downto 0);
  signal offgain_1_3_offset   : std_logic_vector(15 downto 0);
  signal algnd_sync           : std_logic_vector(3 downto 0);
  signal algnd_data           : std_logic_vector(63 downto 0);
  signal cal_trigger          : std_logic;
  signal dac_shift_cnt_l      : std_logic_vector(3 downto 0);
  signal sw_trig_xdom         : std_logic;
  signal sw_trig_demet        : std_logic;
  signal sw_cal_trig          : std_logic;
  signal sel_trig_mode        : std_logic_vector(2 downto 0);
  signal test_data_req        : std_logic;
  signal test_data            : std_logic_vector(63 downto 0);
  signal test_data_vld        : std_logic;
  signal pattern_test         : std_logic;

begin

  -- Synchronize dac_reset to dac_clk_bufr_l domain
  process (dac_reset, dac_clk_bufr_l)
  begin
    if (dac_reset = '1') then
      dac_rst_sreg <= (others => '1');
    elsif (rising_edge(dac_clk_bufr_l)) then
      dac_rst_sreg <= dac_rst_sreg(dac_rst_sreg'high-1 downto 0) & '0';
    end if;
  end process;

  phy_rst <= dac_rst_sreg(dac_rst_sreg'high);

  -- fifo_rst must be set for at least 3 write and read clock cycles
  -- therefore tieing it to dac_run ensures this condition is met
  fifo_rst <= not dac_run;

  -- select either input data or test data
  process (sys_clk)
  begin
    if (rising_edge(sys_clk)) then
      if (srst = '1' or dac_run = '0') then
        selected_wr  <= '0';
        selected_din <= (others => '0');
      elsif (test_en = '1') then
        selected_wr  <= test_data_vld;
        selected_din <= test_data;
      else
        selected_wr  <= din_wr;
        selected_din <= din;
      end if;
    end if;
  end process;

  -- Mux the gain and offset coefficients of the odd numbered samples
  -- to apply DAC-A coefficients when in single channel mode and DAC-B
  -- coefficients when in dual channel mode.
  -- Also force all these coefficients to default values when in pattern
  -- test mode to not get modified values out of the offgain component when
  -- in this test mode which will cause the test to fail.
  offgain_0_2_gain   <= ("01" & x"0000") when (pattern_test = '1') else
                        dac_a_gain;
  offgain_0_2_offset <= x"0000" when (pattern_test = '1') else
                        dac_a_offset;
  offgain_1_3_gain   <= ("01" & x"0000") when (pattern_test = '1') else
                        dac_b_gain when (dac_dual_ch = '1') else
                        dac_a_gain;
  offgain_1_3_offset <= x"0000" when (pattern_test = '1') else
                        dac_b_offset when (dac_dual_ch = '1') else
                        dac_a_offset;

  -- Offset and gain correction
  inst_offgain_0 : ii_offgain
    port map (
      srst                 => srst,
      clk                  => sys_clk,
      gain                 => offgain_0_2_gain,
      offset               => offgain_0_2_offset,
      ce                   => selected_wr,
      din                  => selected_din(15 downto 0),
      data_vld             => offgain_vld,
      dout                 => offgain_dout(15 downto 0)
    );

  inst_offgain_1 : ii_offgain
    port map (
      srst                 => srst,
      clk                  => sys_clk,
      gain                 => offgain_1_3_gain,
      offset               => offgain_1_3_offset,
      ce                   => selected_wr,
      din                  => selected_din(31 downto 16),
      data_vld             => open,
      dout                 => offgain_dout(31 downto 16)
    );

  inst_offgain_2 : ii_offgain
    port map (
      srst                 => srst,
      clk                  => sys_clk,
      gain                 => offgain_0_2_gain,
      offset               => offgain_0_2_offset,
      ce                   => selected_wr,
      din                  => selected_din(47 downto 32),
      data_vld             => open,
      dout                 => offgain_dout(47 downto 32)
    );

  inst_offgain_3 : ii_offgain
    port map (
      srst                 => srst,
      clk                  => sys_clk,
      gain                 => offgain_1_3_gain,
      offset               => offgain_1_3_offset,
      ce                   => selected_wr,
      din                  => selected_din(63 downto 48),
      data_vld             => open,
      dout                 => offgain_dout(63 downto 48)
    );

  -- store corrected data in a fifo
  inst_dac_fifo : afifo_512x64_bram
    port map (
      rst                  => fifo_rst,
      wr_clk               => sys_clk,
      rd_clk               => dac_clk_bufr_l,
      din                  => offgain_dout,
      wr_en                => offgain_vld,
      rd_en                => fifo_rden,
      dout                 => fifo_dout,
      full                 => open,
      empty                => open,
      valid                => fifo_dout_vld,
      underflow            => fifo_underflow,
      prog_full            => fifo_afull
    );

  process (sys_clk)
  begin
    if (rising_edge(sys_clk)) then
      fifo_afull_d <= fifo_afull;
      fifo_rdy_l   <= not fifo_afull_d and dac_run;
    end if;
  end process;

  fifo_rdy <= fifo_rdy_l;

-----------------------------------------------------------------------------
-- FIFO Underflow logic
-----------------------------------------------------------------------------
  -- generate underflow level signal @ dac_clk_bufr_l domain
  process (srst, dac_clk_bufr_l)
  begin
    if (srst = '1') then      -- srst is synchronous to sys_clk domain
      underflow_latch   <= '0';
    elsif (rising_edge(dac_clk_bufr_l)) then
      if (fifo_underflow = '1') then
        assert (false) report "DAC fifo underflow!" severity error;
        underflow_latch <= '1';
      end if;
    end if;
  end process;

  -- Sync underflow latch level signal to sys_clk domain
  -- and generate underflow level signal for alert
  process (sys_clk)
  begin
    if (rising_edge(sys_clk)) then
      if (srst = '1') then
        underflow_latch_xdom  <= '0';
        underflow_latch_demet <= '0';
      else
        underflow_latch_xdom  <= underflow_latch;
        underflow_latch_demet <= underflow_latch_xdom;
      end if;
    end if;
  end process;

  underflow <= underflow_latch_demet;
-----------------------------------------------------------------------------

-----------------------------------------------------------------------------
-- Instantiate ii_trigger
-----------------------------------------------------------------------------
  inst_trigger : ii_trigger
    generic map (
      SAMPLES_PER_CLK      => 1
    )
    port map (
      reset                => phy_rst,
      clk                  => dac_clk_bufr_l,
      ce                   => dac_run,
      ext_sync             => ext_sync,
      sw_trig              => sw_cal_trig,
      trig_mode            => sel_trig_mode,
      frame_size           => window_size,
      decimation_coeff     => (others => '0'),
      decimation_en        => open,
      trigger              => trigger,
      trigger_en           => dac_trigger_en
    );
-----------------------------------------------------------------------------

  -- Toggle ph_en when dac_dll_bypass is set
  process (dac_clk_bufr_l)
  begin
    if (rising_edge(dac_clk_bufr_l)) then
      if (dac_dll_bypass = '1') then
        ph_en <= not ph_en;
      else
        ph_en <= '1';
      end if;
    end if;
  end process;

  fifo_rden <= trigger and ph_en;

  -- fifo data valid generates the sync_out signal
  process (srst, dac_clk_bufr_l)
  begin
    if (srst = '1') then      -- srst is synchronous to sys_clk domain
      fifo_dout_vld_d  <= '0';
      fifo_dout_vld_dd <= '0';
    elsif (rising_edge(dac_clk_bufr_l)) then
      fifo_dout_vld_d  <= fifo_dout_vld;
      fifo_dout_vld_dd <= fifo_dout_vld_d;
    end if;
  end process;

  -- register the fifo output to ease timing
  process (dac_clk_bufr_l)
  begin
    if (rising_edge(dac_clk_bufr_l)) then
      fifo_underflow_d  <= fifo_underflow;
      fifo_underflow_dd <= fifo_underflow_d;
      if (dac_run = '0') then
        fifo_dout_d <= (others => '0');
      elsif (fifo_dout_vld = '1' and fifo_underflow = '0') then
        fifo_dout_d <= fifo_dout;
      end if;
    end if;
  end process;

  -- raw_sync should be set during fifo_dout_vld_d and while
  -- loading the upper words when dac_dll_bypass is asserted
  raw_sync <= (dac_dll_bypass and fifo_dout_vld_dd) or
              fifo_dout_vld_d;

  -- Mux the input to the PHY so that zeros are transmitted whenever
  -- raw_sync deasserts.
  -- Also repeat each sample twice when dac_dll_bypass is asserted
  process (fifo_dout_d, raw_sync, dac_dll_bypass, dac_dual_ch,
           fifo_dout_vld_d, fifo_underflow_d, fifo_underflow_dd)
  begin
    if (raw_sync = '0') then
      raw_data <= (others => '0');
    elsif ((fifo_underflow_dd = '1' and dac_dll_bypass = '1') or
           fifo_underflow_d = '1') then   -- repeat the last sample
      if (dac_dual_ch = '1') then
        if (dac_dll_bypass = '1') then
          raw_data <= fifo_dout_d(63 downto 48) & fifo_dout_d(63 downto 48) &
                      fifo_dout_d(47 downto 32) & fifo_dout_d(47 downto 32);
        else
          raw_data <= (fifo_dout_d(63 downto 32) & fifo_dout_d(63 downto 32));
        end if;
      else
        raw_data <= (fifo_dout_d(63 downto 48) & fifo_dout_d(63 downto 48) &
                    fifo_dout_d(63 downto 48) & fifo_dout_d(63 downto 48));
      end if;
    elsif (dac_dll_bypass = '0') then     -- load 4 samples on every clock
      raw_data <= fifo_dout_d;
    else                                  -- repeat each word twice
      if (fifo_dout_vld_d = '1') then     -- repeat and load the lower words
        raw_data <= fifo_dout_d(31 downto 16) & fifo_dout_d(31 downto 16) &
                    fifo_dout_d(15 downto 0) & fifo_dout_d(15 downto 0);
      else                                -- repeat and load the upper words
        raw_data <= fifo_dout_d(63 downto 48) & fifo_dout_d(63 downto 48) &
                    fifo_dout_d(47 downto 32) & fifo_dout_d(47 downto 32);
      end if;
    end if;
  end process;
  -----------------------------------------------------------------------------

-----------------------------------------------------------------------------
-- dac_trig_alrt alert logic
-----------------------------------------------------------------------------
  -- detect a rising edge on trigger @dac_clk_bufr_l domain
  process (dac_clk_bufr_l)
  begin
    if (rising_edge(dac_clk_bufr_l)) then
      trigger_d <= trigger;
    end if;
  end process;

  trigger_re <= not trigger_d and trigger;

  -- generate trigger latch level signal @dac_clk_bufr_l domain
  -- on the first rising edge of trigger after a reset
  process (srst, dac_clk_bufr_l)
  begin
    if (srst = '1') then      -- srst is synchronous to sys_clk domain
      trigger_latch   <= '0';
    elsif (rising_edge(dac_clk_bufr_l)) then
      if (trigger_re = '1') then
        trigger_latch <= '1';
      end if;
    end if;
  end process;

  -- Sync trigger_latch level signal to sys_clk domain
  -- and generate dac_trig_alrt level signal for alert
  process (sys_clk)
  begin
    if (rising_edge(sys_clk)) then
      if (srst = '1') then
        trigger_latch_xdom  <= '0';
        trigger_latch_demet <= '0';
      else
        trigger_latch_xdom  <= trigger_latch;
        trigger_latch_demet <= trigger_latch_xdom;
      end if;
    end if;
  end process;

  dac_trig_alrt <= trigger_latch_demet;
-----------------------------------------------------------------------------

-----------------------------------------------------------------------------
-- Instantiate ii_dac_bitslip
-----------------------------------------------------------------------------
  -- Latch the phase of the dac clock on the rising edge of trigger
  process (dac_clk_bufr_l)
  begin
    if (rising_edge(dac_clk_bufr_l)) then
      if (trigger_re = '1') then
        trig_clk_phase <= ph_en;
      end if;
    end if;
  end process;

  dac_bitslip_inst : ii_dac_bitslip
    port map (
      -- clock
      dac_clk_bufr         => dac_clk_bufr_l,

      -- control
      trig_clk_phase       => trig_clk_phase,
      dac_dual_ch          => dac_dual_ch,
      dac_dll_bypass       => dac_dll_bypass,
      dac_shift_cnt        => dac_shift_cnt_l,
      ext_sync_phase       => ext_sync_phase,

      -- raw DAC data
      raw_sync             => raw_sync,
      raw_data             => raw_data,

      -- aligned DAC data
      algnd_sync           => algnd_sync,
      algnd_data           => algnd_data
    );
-----------------------------------------------------------------------------

-----------------------------------------------------------------------------
-- Instantiate ii_dac5682z_phy
-----------------------------------------------------------------------------
  dac5682z_phy_inst : ii_dac5682z_phy
    port map (
      phy_rst              => phy_rst,
      idelayctrl_rst       => idelayctrl_rst,
      ref_clk200           => ref_clk200,
      dac_clk_bufio        => dac_clk_bufio_l,
      dac_clk_bufr         => dac_clk_bufr_l,
      dac_dll_bypass       => dac_dll_bypass,

      -- Parallel data and output enable
      sync_in              => algnd_sync,
      data_in              => algnd_data,

      -- DAC interface signals
      dac_clk_in_p         => dac_clk_in_p,
      dac_clk_in_n         => dac_clk_in_n,
      dac_clk_out_p        => dac_clk_out_p,
      dac_clk_out_n        => dac_clk_out_n,
      sync_out_p           => sync_out_p,
      sync_out_n           => sync_out_n,
      sync2_out_p          => sync2_out_p,
      sync2_out_n          => sync2_out_n,
      data_out_p           => data_out_p,
      data_out_n           => data_out_n
    );

  dac_clk_bufio <= dac_clk_bufio_l;
  dac_clk_bufr  <= dac_clk_bufr_l;
-----------------------------------------------------------------------------

-----------------------------------------------------------------------------
-- Instantiate ii_dac_lat_cal
-----------------------------------------------------------------------------
  lat_cal_inst : ii_dac_lat_cal
    port map (
      -- Reset and clocks
      dac_reset            => dac_reset,
      fs_clk               => dac_clk_bufio_l,
      fs_clkdiv2           => dac_clk_bufr_l,

      -- Controls
      dac_cal_en           => dac_cal_en,
      dac_run              => dac_run,
      dac_dual_ch          => dac_dual_ch,
      dac_dll_bypass       => dac_dll_bypass,

      -- DAC output digitizer interface
      dac_dig_p            => dac_dig_p,
      dac_dig_n            => dac_dig_n,

      -- Outputs
      cal_trigger          => cal_trigger,
      dac_cal0_done        => dac_cal0_done,
      dac_cal1_done        => dac_cal1_done,
      dac_iodly_cnt        => dac_iodly_cnt,
      dac_shift_cnt        => dac_shift_cnt_l
    );

  dac_shift_cnt <= dac_shift_cnt_l;

  -- Sync the software trigger to dac_clk_bufr_l domain and
  -- logical OR it with the latency calibration module's
  -- trigger output. Connect the resulting trigger to the software
  -- trigger port of the trigger module
  process (dac_clk_bufr_l)
  begin
    if (rising_edge(dac_clk_bufr_l)) then
      sw_trig_xdom  <= sw_trig;
      sw_trig_demet <= sw_trig_xdom;
      sw_cal_trig   <= (sw_trig_demet and not dac_cal_en) or cal_trigger;
    end if;
  end process;

  -- Override the trigger mode signal when running the DAC calibration
  process (sys_clk)
  begin
    if (rising_edge(sys_clk)) then
      if (dac_cal_en = '1') then
        sel_trig_mode <= (others => '0');
      else
        sel_trig_mode <= trigger_mode;
      end if;
    end if;
  end process;
-----------------------------------------------------------------------------

-----------------------------------------------------------------------------
-- Instantiate DAC test data generator
-----------------------------------------------------------------------------
  -- request test data from the test generator
  process (sys_clk)
  begin
    if (rising_edge(sys_clk)) then
      if (srst = '1') then
        test_data_req <= '0';
      else
        test_data_req <= fifo_rdy_l and test_en;
      end if;
    end if;
  end process;

  inst_dac_test_gen : ii_dac_test_gen
  port map (
    -- Reset and clock
    srst            => srst,
    sys_clk         => sys_clk,

    -- Control
    test_en         => test_en,
    test_mode       => test_mode,
    phase_inc_wr    => phase_inc_wr,
    phase_inc       => phase_inc,

    -- Data
    test_data_req   => test_data_req,
    dout            => test_data,
    valid           => test_data_vld,
    pattern_test    => pattern_test
  );
-----------------------------------------------------------------------------

end arch;
