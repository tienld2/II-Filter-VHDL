-------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   15:34:34 09/05/2013
-- Design Name:   
-- Module Name:   /home/nick/polyDecimDemodFilter/polyDecimDemodFilter_Top_tb.vhd
-- Project Name:  polyDecimDemodFilter
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: polyDecimDemodFilter_Top
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
use IEEE.std_logic_misc.all;
use IEEE.std_logic_unsigned.all;

library ieee_proposed;
use ieee_proposed.fixed_float_types.all;
use ieee_proposed.fixed_pkg.all;

 
ENTITY polyDecimDemodFilter_Top_tb IS
END polyDecimDemodFilter_Top_tb;
 
ARCHITECTURE behavior OF polyDecimDemodFilter_Top_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT polyDecimDemodFilter_Top
    PORT(
         clk : IN  std_logic;
         clk_enable : IN  std_logic;
         max_count : IN unsigned(3 downto 0);
         rst : IN  std_logic;
         tValidIn_Array : IN  std_logic_vector(15 downto 0);
         runSignals : IN  std_logic_vector(15 downto 0);
         numTaps : IN  std_logic_vector(4 downto 0);
         decimFactor : IN  real;
         reloadCoefData : IN  std_logic_vector(15 downto 0);
         phaseInc : IN  std_logic_vector(15 downto 0);
         inputSignal : IN  std_logic_vector(15 downto 0);
         -- -------------------------------------------------
         -- temporary signals -------------------------------
         datatoDemodTop : out std_logic_vector(15 downto 0) ;
         dataOutFromDemodRe : out std_logic_vector(31 downto 0) ;
         dataOutFromDemodIm  : out std_logic_vector(31 downto 0) ;
         -- temporary signals -------------------------------
         -- -------------------------------------------------
         outputDataRe : OUT  std_logic_vector(15 downto 0);
         outputDataIm : OUT  std_logic_vector(15 downto 0)
        );
    END COMPONENT;


   function cast_to_signed_int16(signal slv: std_logic_vector) return signed is
   begin
     return to_signed(to_integer(signed(slv)),16);
   end cast_to_signed_int16;

    
   --Inputs
   signal clk : std_logic := '0';
   signal clk_enable : std_logic := '0';
   signal clk_div : std_logic := '0';                         --   (samplingFreq / decimFactor) / 2
   signal max_count : unsigned(3 downto 0) := b"0001";   --   (100 MHz      / 4          ) / 2 = 12500000 
   signal rst : std_logic := '0';
   signal tValidIn_Array : std_logic_vector(15 downto 0) := (others => '0');
   signal runSignals : std_logic_vector(15 downto 0) := (others => '0');
   signal numTaps : std_logic_vector(4 downto 0) := (others => '0');
   signal decimFactor : real := 4.0;
   signal reloadCoefData : std_logic_vector(15 downto 0) := (others => '0');
   signal phaseInc : std_logic_vector(15 downto 0) := (others => '0');
   signal inputSignal : std_logic_vector(15 downto 0) := (others => '0');
   -- -------------------------------------------------
   -- temporary signals -------------------------------
   signal datatoDemodTop : std_logic_vector(15 downto 0) := (others => '0');
   signal dataOutFromDemodRe : std_logic_vector(31 downto 0) := (others => '0');
   signal dataOutFromDemodIm  : std_logic_vector(31 downto 0) := (others => '0');
   -- temporary signals -------------------------------
   -- -------------------------------------------------


  -- Constants
  constant inputSize : integer := 4095;

 	--Outputs
   signal outputDataRe : std_logic_vector(15 downto 0);
   signal outputDataIm : std_logic_vector(15 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
   constant clk_enable_period : time := 10 ns;

    -- clock divided clock:
    signal clk_div_counter : integer := 0;
    signal clk_div_temp : std_logic := '1';


  type input_array is array (0 to inputSize) of std_logic_vector(15 downto 0) ;
signal myCosine : input_array :=(x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000");

BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: polyDecimDemodFilter_Top PORT MAP (
          clk => clk,
          clk_enable => clk_enable,
          max_count => max_count,
          rst => rst,
          tValidIn_Array => tValidIn_Array,
          runSignals => runSignals,
          numTaps => numTaps,
          decimFactor => decimFactor,
          reloadCoefData => reloadCoefData,
          phaseInc => phaseInc,
          inputSignal => inputSignal,
          -- -------------------------------------------------
          -- temporary signals -------------------------------
          datatoDemodTop => datatoDemodTop,
          dataOutFromDemodRe => dataOutFromDemodRe,
          dataOutFromDemodIm => dataOutFromDemodIm,
          -- temporary signals -------------------------------
          -- -------------------------------------------------
          outputDataRe => outputDataRe,
          outputDataIm => outputDataIm
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 
   clk_enable_process :process
   begin
		clk_enable <= '0';
		wait for clk_enable_period/2;
		clk_enable <= '1';
		wait for clk_enable_period/2;
   end process;


   -- ------------------------------------------------------------------------------------------------------
   --                                       temporary signals 
   -- ------------------------------------------------------------------------------------------------------
   output_filedatatoDemodTop : entity work.file_writer 
   generic map( 
     dataWidth => 16,
     wordWidth => 1,
     -- dataFrac => 15,
     fileName => "/home/nick/polyDecimDemodFilter/dataFromFIRFilteroutput10MHz.dat"
   )
   port map( 
     reset => rst,
     clk => clk_div,
     enable => tValidIn_Array(0),
     data => datatoDemodTop,
     data_valid => tValidIn_Array(0)
   );

   output_filedataDemodReoutput : entity work.file_writer 
   generic map( 
     dataWidth => 16,
     wordWidth => 1,
     -- dataFrac => 15,
     fileName => "/home/nick/polyDecimDemodFilter/dataDemodReoutput10MHz.dat"
   )
   port map( 
     reset => rst,
     clk => clk_div,
     enable => tValidIn_Array(0),
     data => dataOutFromDemodRe(31 downto 16),-- to_slv(to_SFix(dataOutFromDemodRe(31 downto 16),16,15)),
     data_valid => tValidIn_Array(0)
   );

   output_filedataDemodImoutput : entity work.file_writer 
   generic map( 
     dataWidth => 16,
     wordWidth => 1,
     -- dataFrac => 15,
     fileName => "/home/nick/polyDecimDemodFilter/dataDemodImoutput10MHz.dat"
   )
   port map( 
     reset => rst,
     clk => clk_div,
     enable => tValidIn_Array(0),
     data => dataOutFromDemodIm(31 downto 16),--to_slv(to_SFix(dataOutFromDemodIm(31 downto 16),16,15)),
     data_valid => tValidIn_Array(0)
   );
   -- ------------------------------------------------------------------------------------------------------
   -- ------------------------------------------------------------------------------------------------------



   -- clk for file writer from iir filters:
   my_clk_div : entity work.clk_div_top
    port map(
      max_count => max_count,
      clk_in => clk,
      rst => rst,
      clk_out => clk_div
    ) ;

  output_fileCos : entity work.file_writer 
  generic map( 
    dataWidth => 16,
    wordWidth => 1,
    -- dataFrac => 15,
    fileName => "/home/nick/polyDecimDemodFilter/cosoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk_div,
    enable => tValidIn_Array(0),
    data => inputSignal,
    data_valid => tValidIn_Array(0)
  );


  -- ------------------------------------------------------------------------------------------------------
  --                        plotted with plotChannelizer.py
  -- ------------------------------------------------------------------------------------------------------

  output_fileRe : entity work.file_writer 
  generic map( 
    dataWidth => 16,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/polyDecimDemodFilter/polyDecimDemodFilterReoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk_div,
    enable => '1',
    data => outputDataRe,
    data_valid => '1'
  );

  output_fileIm : entity work.file_writer 
  generic map( 
    dataWidth => 16,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/polyDecimDemodFilter/polyDecimDemodFilterImoutput10MHz.dat"
  )
  port map( 
    reset => rst,
    clk => clk_div,
    enable => '1',
    data => outputDataIm,
    data_valid => '1'
  );

  -- ------------------------------------------------------------------------------------------------------
  -- ------------------------------------------------------------------------------------------------------



   -- Stimulus process
   stim_proc: process
   begin		

      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;

      -- insert, stimulus here 
      -- pulse the reset line:
      rst <= '1'; wait until (rising_edge(clk));
      wait for clk_period*4;
      rst <= '0'; wait until (rising_edge(clk));
      report "System reset with global signal rst.\n";


      -- feed data into polyDecimator, start filtering:
      tValidIn_Array(0) <= '1'; wait until (rising_edge(clk));
      runSignals(0) <= '1'; wait until (rising_edge(clk));
      report "polyDecimator triggered, transmitting data to filter now...\n";

      tValidIn_Array(1) <= '1';
						phaseInc <= x"147A"; wait until (rising_edge(clk));						
            -- phaseInc <= x"0000"; wait until (rising_edge(clk));           

      for i in 0 to inputSize loop
        inputSignal <= myCosine(i); wait until (rising_edge(clk)); 
      end loop;



      -- initiate demodulator when signal available from filter, set phaseInc:
      

      report "Setting phaseInc to 0x0CCC, initiating demodulator...\n";

      report "Finished processing.";

      wait;
   end process;

END;
