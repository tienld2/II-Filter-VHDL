-------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   15:34:34 09/05/2013
-- Design Name:   
-- Module Name:   /home/nick/polyDecimDemodFilter2/polyDecimDemodFilter2_Top_tb.vhd
-- Project Name:  polyDecimDemodFilter2
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: polyDecimDemodFilter2_Top
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_textio.all;

library STD;
use std.textio.all;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
-- USE ieee.numeric_std.ALL;
 
use work.mappings.all;
use work.parameters.all;


ENTITY polyDecimDemodFilter2_Top_tb IS
END polyDecimDemodFilter2_Top_tb;
 
ARCHITECTURE behavior OF polyDecimDemodFilter2_Top_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT polyDecimDemodFilter2_Top
    PORT(
      clk1                  : in    std_logic;
      hi_in                 : in    std_logic_vector(7 downto 0);
      hi_out                : out   std_logic_vector(1 downto 0);
      hi_inout              : inout std_logic_vector(15 downto 0);
      hi_muxsel             : out   std_logic;
      i2c_sda               : out   std_logic;
      i2c_scl               : out   std_logic;
      led                   : out   std_logic_vector(7 downto 0);
      -- -------------------------------------------------
      -- temporary signals -------------------------------
      -- acc_padRe             : out std_logic_vector(49 downto 0); 
      -- acc_padIm             : out std_logic_vector(49 downto 0);
      inputSignalBis        : out std_logic_vector(15 downto 0);
      datatoDemodTop        : out std_logic_vector(19 downto 0);
      dataOutFromDemodRe    : out std_logic_vector(35 downto 0);
      dataOutFromDemodIm    : out std_logic_vector(35 downto 0);
      mulOutput             : out std_logic_vector(79 downto 0);
      blockRamOutput        : out std_logic_vector(31 downto 0);
      iirFilterTmp          : out std_logic_vector(39 downto 0) 
      -- temporary signals -------------------------------
      -- -------------------------------------------------

  );
    END COMPONENT;

  --Inputs
  signal wireInLines        : std_logic_vector(15 downto 0) := (others => '0');
  signal ti_clk             : std_logic;
  signal slow_clk           : std_logic_vector(15 downto 0) ;
  signal clk_enable         : std_logic := '0';     -- (samplingFreq / decimFactor) / 2
  signal clk_div            : std_logic := '0';     -- (    100 MHz  / 4 ) / 2 = 12500000 
  signal max_count          : natural := 1;         
  signal tValidIn_Array     : std_logic_vector(15 downto 0) := (others => '0');
  signal runSignals         : std_logic_vector(15 downto 0) := (others => '0');
  signal reloadFIRCoefData  : std_logic_vector(15 downto 0) := (others => '0');
  signal phaseInc           : std_logic_vector(15 downto 0) := (others => '0');
  signal inputSignal        : std_logic_vector(15 downto 0) := (others => '0');
  signal inputSignalBis     : std_logic_vector(15 downto 0) := (others => '0');
  signal windowCoef         : std_logic_vector(31 downto 0);
  signal trigger_array      : std_logic_vector(4 downto 0);
  signal decimFactor        : natural := 4;

  --Inputs
  signal hi_in              : std_logic_vector(7 downto 0) := (others => '0');
  signal clk1               : std_logic := '0';
  signal ok1                : std_logic_vector(30 downto 0);
  signal ok2                : std_logic_vector(16 downto 0);
  signal ok2s               : std_logic_vector(17*10-1 downto 0);
  

  --BiDirs
  signal hi_inout           : std_logic_vector(15 downto 0);
  signal hi_aa              : std_logic;

  --Outputs
  signal hi_out             : std_logic_vector(1 downto 0);
  signal hi_muxsel          : std_logic;
  signal i2c_sda            : std_logic;
  signal i2c_scl            : std_logic;
  signal led                : std_logic_vector(7 downto 0);

  signal hi_clk             : std_logic;
  signal hi_dataout         : std_logic_vector(15 downto 0) := x"0000";

  -- Clock periods
  constant clk1_period      : time := 10 ns;      -- 100 MHz clk period
  constant tCK              : time := 10.417 ns;  -- half period for 48 MHz
  constant clk_en_period    : time := 10 ns;
  constant clk_div_period   : time := 40 ns;

  -- Constants
  constant inputSize        : integer := 4095;
  constant windowSize       : integer := 1023;

  --Outputs
  signal outputDataRe       : std_logic_vector(19 downto 0);
  signal outputDataIm       : std_logic_vector(19 downto 0);
  signal acc                : std_logic_vector(99 downto 0);

  -- -------------------------------------------------  
  -- temporary signals -------------------------------
  signal acc_padRe          : std_logic_vector(49 downto 0) := (others => '0');
  signal acc_padIm          : std_logic_vector(49 downto 0) := (others => '0');
  signal datatoDemodTop     : std_logic_vector(19 downto 0) := (others => '0');
  signal dataOutFromDemodRe : std_logic_vector(35 downto 0) := (others => '0');
  signal dataOutFromDemodIm : std_logic_vector(35 downto 0) := (others => '0');
  signal mulOutput          : std_logic_vector(79 downto 0);
  signal blockRamOutput     : std_logic_vector(31 downto 0);
  signal iirFilterTmp       : std_logic_vector(39 downto 0);
  -- temporary signals -------------------------------
  -- -------------------------------------------------

  -- signals to file writer
  signal acc_padRe2         : std_logic_vector(63 downto 0) := (others => '0');
  signal acc_padIm2         : std_logic_vector(63 downto 0) := (others => '0');
  signal padding            : std_logic_vector(13 downto 0) := (others => '0');
  signal accReLSB, accImLSB : std_logic_vector(31 downto 0);


  -- inputSize, windowSize = total lengths of input and window coefficients
  type input_array is array (0 to inputSize) of std_logic_vector(15 downto 0);
  type input_array32 is array (0 to windowSize) of std_logic_vector(31 downto 0);
  signal myCosine : input_array := (x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"E805",x"F7F7",x"0809",x"17FB",x"278D",x"367F",x"4495",x"5196",x"5D4E",x"678D",x"7029",x"7701",x"7BF9",x"7EFC",x"7FFF",x"7EFC",x"7BF9",x"7701",x"7029",x"678D",x"5D4E",x"5196",x"4495",x"367F",x"278D",x"17FB",x"0809",x"F7F7",x"E805",x"D873",x"C981",x"BB6B",x"AE6A",x"A2B2",x"9873",x"8FD7",x"88FF",x"8407",x"8104",x"8001",x"8104",x"8407",x"88FF",x"8FD7",x"9873",x"A2B2",x"AE6A",x"BB6B",x"C981",x"D873",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"8246",x"8042",x"8042",x"8246",x"8645",x"8C30",x"93EE",x"9D61",x"A862",x"B4C5",x"C257",x"D0E2",x"E02C",x"EFF6",x"0000",x"100A",x"1FD4",x"2F1E",x"3DA9",x"4B3B",x"579E",x"629F",x"6C12",x"73D0",x"79BB",x"7DBA",x"7FBE",x"7FBE",x"7DBA",x"79BB",x"73D0",x"6C12",x"629F",x"579E",x"4B3B",x"3DA9",x"2F1E",x"1FD4",x"100A",x"0000",x"EFF6",x"E02C",x"D0E2",x"C257",x"B4C5",x"A862",x"9D61",x"93EE",x"8C30",x"8645",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000");
   -- signal myCoef : input_array32 :=(x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"0000FFFF",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");
   signal myCoef : input_array32 := (others => x"00007fff");

BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: polyDecimDemodFilter2_Top PORT MAP (
      clk1   => clk1,
      hi_in    => hi_in,
      hi_out   => hi_out,
      hi_inout => hi_inout,
      hi_muxsel=> hi_muxsel,
      i2c_sda  => i2c_sda,
      i2c_scl  => i2c_scl,
      led      => led,
  -- -------------------------------------------------
  -- temporary signals -------------------------------
  -- acc_padRe =>  acc_padRe,
  -- acc_padIm   => acc_padIm ,
  inputSignalBis => inputSignalBis,
  datatoDemodTop => datatoDemodTop,
  dataOutFromDemodRe => dataOutFromDemodRe,
  dataOutFromDemodIm  => dataOutFromDemodIm ,
  mulOutput => mulOutput,
  blockRamOutput => blockRamOutput,
  iirFilterTmp => iirFilterTmp
  -- temporary signals -------------------------------
  -- -------------------------------------------------
  );

 
  hi_in(0) <= hi_clk;
  hi_inout <= hi_dataout when (hi_in(1) = '1') else (others => 'Z');
 

  -- concatenate 50 & 50 = 100 bits
  -- acc <= acc_padIm & acc_padRe;

 
  -- Clock Generation Process
  hi_clk_gen : process is
  begin
    hi_clk <= '0';
    wait for tCk;
    hi_clk <= '1'; 
    wait for tCk; 
  end process hi_clk_gen;

  -- 100 MHz clock, 50% duty cycle:
  clk_process :process
  begin
    clk1 <= '0';
    wait for clk1_period/2;
    clk1 <= '1';
    wait for clk1_period/2;
  end process;

 
   clk_enable_process :process
   begin
    clk_enable <= '0';
    wait for clk_en_period/2;
    clk_enable <= '1';
    wait for clk_en_period/2;
   end process;

   -- clk for file writer from iir filters:
   my_clk_div : entity work.clk_div_top
    port map(
      max_count => max_count,
      clk_in => clk1,
      rst => wireInLines(0),
      clk_out => clk_div
    );


-- ----------------------------------------------------------------------------------------------
--                              File Writer Block
-- ----------------------------------------------------------------------------------------------

-- -------------------------------------- 
--        Input Signal File Writer
-- --------------------------------------
output_fileCos : entity work.file_writer 
  generic map( 
    dataWidth => 16,
    wordWidth => 1,
    -- dataFrac => 15,
    fileName => "/home/nick/polyDecimDemodFilter2/cosoutput10MHz.dat"
  )
  port map( 
    reset => wireInLines(0),
    clk => clk1,
    enable => wireInLines(2),
    data => inputSignalBis,
    data_valid => wireInLines(2)
  );

-- -------------------------------------- 
--   Polyphase FIRFilter File Writer
-- --------------------------------------
output_filedatatoDemodTop : entity work.file_writer 
  generic map( 
    dataWidth => 20,
    wordWidth => 1,
    -- dataFrac => 15,
    fileName => "/home/nick/polyDecimDemodFilter2/dataFromFIRFilteroutput10MHz.dat"
  )
  port map( 
    reset => wireInLines(0),
    clk => clk_div,
    enable => wireInLines(3),
    data => datatoDemodTop,
    data_valid => wireInLines(3)
  );

-- -------------------------------------- 
--        Demodulator File Writers
-- --------------------------------------
output_filedataDemodReoutput : entity work.file_writer 
  generic map( 
     dataWidth => 20,
     wordWidth => 1,
     -- dataFrac => 15,
     fileName => "/home/nick/polyDecimDemodFilter2/dataDemodReoutput10MHz.dat"
  )
  port map( 
     reset => wireInLines(0),
     clk => clk_div,
     enable => wireInLines(3),
     data => dataOutFromDemodRe(30 downto 11),
     data_valid => wireInLines(3)
  );
output_filedataDemodImoutput : entity work.file_writer 
  generic map( 
     dataWidth => 20,
     wordWidth => 1,
     -- dataFrac => 15,
     fileName => "/home/nick/polyDecimDemodFilter2/dataDemodImoutput10MHz.dat"
  )
  port map( 
     reset => wireInLines(0),
     clk => clk_div,
     enable => wireInLines(3),
     data => dataOutFromDemodIm(30 downto 11),
     data_valid => wireInLines(3)
  );


-- -------------------------------------- 
--        IIRFilter File Writers
-- --------------------------------------
output_fileiirreal : entity work.file_writer 
  generic map( 
    dataWidth => 20,
    wordWidth => 1,
    -- dataFrac => 15,
    fileName => "/home/nick/polyDecimDemodFilter2/dataIIRFilterReoutput10MHz.dat"
  )
  port map( 
    reset => wireInLines(0),
    clk => clk_div,
    enable => wireInLines(2),
    data => iirFilterTmp(19 downto 0),
    data_valid => wireInLines(2)
  );
output_fileiirimag : entity work.file_writer 
  generic map( 
    dataWidth => 20,
    wordWidth => 1,
    -- dataFrac => 15,
    fileName => "/home/nick/polyDecimDemodFilter2/dataIIRFilterImoutput10MHz.dat"
  )
  port map( 
    reset => wireInLines(0),
    clk => clk_div,
    enable => wireInLines(2),
    data => iirFilterTmp(39 downto 20),
    data_valid => wireInLines(2)
  );

-- -------------------------------------- 
--        Window Function File Writer
-- --------------------------------------
output_fileWindow : entity work.file_writer 
  generic map( 
    dataWidth => 32,
    wordWidth => 1,
    -- dataFrac => 15,
    fileName => "/home/nick/polyDecimDemodFilter2/dataMULwindowoutput10MHz.dat"
  )
  port map( 
    reset => wireInLines(0),
    clk => clk_div,
    enable => wireInLines(2),
    data => windowCoef,
    data_valid => wireInLines(2)
  );

-- -------------------------------------- 
--        MUL File Writers
-- --------------------------------------
output_filemulRe : entity work.file_writer 
  generic map( 
    dataWidth => 36,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/polyDecimDemodFilter2/dataMULReoutput10MHz.dat"
  )
  port map( 
    reset => wireInLines(0),
    clk => clk_div,
    enable => wireInLines(2),
    data => mulOutput(35 downto 0),
    data_valid => wireInLines(2)
  );
output_filemulIm : entity work.file_writer 
  generic map( 
    dataWidth => 36,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/polyDecimDemodFilter2/dataMULImoutput10MHz.dat"
  )
  port map( 
    reset => wireInLines(0),
    clk => clk_div,
    enable => wireInLines(2),
    data => mulOutput(75 downto 40),
    data_valid => wireInLines(2)
  );

-- -------------------------------------- 
--        Output Signal File Writers
-- --------------------------------------

-- Bottom 32 bits of outputRe
output_filemacReLSB : entity work.file_writer 
  generic map( 
    dataWidth => 32,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/polyDecimDemodFilter2/polyDecimDemodFilter2ReLSBoutput10MHz.dat"
  )
  port map( 
    reset => wireInLines(0),
    clk => hi_clk,
    enable => wireInLines(2),
    data => acc(31 downto 0),
    data_valid => wireInLines(2)
  );

-- Bottom 32 bits of outputIm
output_filemacImLSB : entity work.file_writer 
  generic map( 
    dataWidth => 32,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/polyDecimDemodFilter2/polyDecimDemodFilter2ImLSBoutput10MHz.dat"
  )
  port map( 
    reset => wireInLines(0),
    clk => hi_clk,
    enable => wireInLines(2),
    data => acc(81 downto 50),
    data_valid => wireInLines(2)
  );

-- Top 18 bits of outputRe
output_filemacReMSB : entity work.file_writer 
  generic map( 
    dataWidth => 18,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/polyDecimDemodFilter2/polyDecimDemodFilter2ReMSBoutput10MHz.dat"
  )
  port map( 
    reset => wireInLines(0),
    clk => hi_clk,
    enable => wireInLines(2),
    data => acc(49 downto 32),
    data_valid => wireInLines(2)
  );

-- Top 18 bits of outputIm
output_filemacImMSB : entity work.file_writer 
  generic map( 
    dataWidth => 18,
    wordWidth => 1,
    -- dataFrac => 10,
    fileName => "/home/nick/polyDecimDemodFilter2/polyDecimDemodFilter2ImMSBoutput10MHz.dat"
  )
  port map( 
    reset => wireInLines(0),
    clk => hi_clk,
    enable => wireInLines(2),
    data => acc(99 downto 82),
    data_valid => wireInLines(2)
  );


-- ----------------------------------------------------------------------------------------------
--                          End of File Writer Block 
-- ----------------------------------------------------------------------------------------------


  --------------------------------------------------------------------------
  -- Begin Simulation Process 
  --------------------------------------------------------------------------
  sim_process : process is

  --<<<<<<<<<<<<<<<<<<< OKHOSTCALLS START PASTE HERE >>>>>>>>>>>>>>>>>>>>-- 
  
-- User defined data for pipe procedures
    -----------------------------------------------------------------------
    variable BlockDelayStates : integer := 5;  -- REQUIRED: # of clocks between blocks of pipe data
    variable ReadyCheckDelay  : integer := 5;  -- REQUIRED: # of clocks before block transfer before
                                               --    host interface checks for ready (0-255)
    variable PostReadyDelay   : integer := 5;  -- REQUIRED: # of clocks after ready is asserted and
                                               --    check that the block transfer begins (0-255)
    variable pipeInSize       : integer := 1024; 
    variable pipeOutSize      : integer := 1024;
  
    -- If you require multiple pipe arrays, you may create more arrays here
    -- duplicate the desired pipe procedures as required, change the names
    -- of the duplicated procedure to a unique identifiers, and alter the
    -- pipe array in that procedure to your newly generated arrays here.
    type PIPEIN_ARRAY is array (0 to pipeInSize - 1) of std_logic_vector(7 downto 0);
    variable pipeIn   : PIPEIN_ARRAY;
  
    type PIPEOUT_ARRAY is array (0 to pipeOutSize - 1) of std_logic_vector(7 downto 0);
    variable pipeOut  : PIPEOUT_ARRAY;
  
    -----------------------------------------------------------------------
    -- Required data for procedures and functions
    -----------------------------------------------------------------------
    type STD_ARRAY is array (0 to 31) of std_logic_vector(15 downto 0);
    variable WireIns, WireOuts, Triggered  :  STD_ARRAY;
  
    constant DNOP                   : std_logic_vector(3 downto 0) := x"0";
    constant DReset                 : std_logic_vector(3 downto 0) := x"1";
    constant DUpdateWireIns         : std_logic_vector(3 downto 0) := x"3";
    constant DUpdateWireOuts        : std_logic_vector(3 downto 0) := x"5";
    constant DActivateTriggerIn     : std_logic_vector(3 downto 0) := x"6";
    constant DUpdateTriggerOuts     : std_logic_vector(3 downto 0) := x"7";
    constant DWriteToPipeIn         : std_logic_vector(3 downto 0) := x"9";
    constant DReadFromPipeOut       : std_logic_vector(3 downto 0) := x"a";
    constant DWriteToBlockPipeIn    : std_logic_vector(3 downto 0) := x"b";
    constant DReadFromBlockPipeOut  : std_logic_vector(3 downto 0) := x"c";
  
    -----------------------------------------------------------------------
    -- FrontPanelReset
    -----------------------------------------------------------------------
    procedure FrontPanelReset is
      variable i : integer := 0;
    begin
        for i in 31 downto 0 loop
          WireIns(i) := (others => '0');
          WireOuts(i) := (others => '0');
          Triggered(i) := (others => '0');
        end loop;
  
        wait until (rising_edge(hi_clk)); hi_in(7 downto 4) <= DReset;
        wait until (rising_edge(hi_clk)); hi_in(7 downto 4) <= DNOP;
        wait until (hi_out(0) = '0');
    end procedure FrontPanelReset;
  
    -----------------------------------------------------------------------
    -- SetWireInValue
    -----------------------------------------------------------------------
    procedure SetWireInValue (
      ep   : in  std_logic_vector(7 downto 0);
      val  : in  std_logic_vector(15 downto 0);
      mask : in  std_logic_vector(15 downto 0)) is
      
      variable tmp_slv16 :     std_logic_vector(15 downto 0);
      variable tmpI      :     integer;
    begin
      tmpI := CONV_INTEGER(ep);
      tmp_slv16 := WireIns(tmpI) and (not mask);
      WireIns(tmpI) := (tmp_slv16 or (val and mask));
    end procedure SetWireInValue;
  
    -----------------------------------------------------------------------
    -- GetWireOutValue
    -----------------------------------------------------------------------
    impure function GetWireOutValue (
      ep : std_logic_vector) return std_logic_vector is
      
      variable tmp_slv16 : std_logic_vector(15 downto 0);
      variable tmpI      : integer;
    begin
      tmpI := CONV_INTEGER(ep);
      tmp_slv16 := WireOuts(tmpI - 16#20#);
      return (tmp_slv16);
    end GetWireOutValue;
  
    -----------------------------------------------------------------------
    -- IsTriggered
    -----------------------------------------------------------------------
    impure function IsTriggered (
      ep   : std_logic_vector;
      mask : std_logic_vector(15 downto 0)) return BOOLEAN is
      
      variable tmp_slv16   : std_logic_vector(15 downto 0);
      variable tmpI        : integer;
      variable msg_line    : line;
    begin
      tmpI := CONV_INTEGER(ep);
      tmp_slv16 := (Triggered(tmpI - 16#60#) and mask);
  
      if (tmp_slv16 >= 0) then
        if (tmp_slv16 = 0) then
          return FALSE;
        else
          return TRUE;
        end if;
      else
        write(msg_line, STRING'("***FRONTPANEL ERROR: IsTriggered mask 0x"));
        hwrite(msg_line, mask);
        write(msg_line, STRING'(" covers unused Triggers"));
        writeline(output, msg_line);
        return FALSE;        
      end if;     
    end IsTriggered;
  
    -----------------------------------------------------------------------
    -- UpdateWireIns
    -----------------------------------------------------------------------
    procedure UpdateWireIns is
      variable i : integer := 0;
    begin
      wait until (rising_edge(hi_clk)); hi_in(7 downto 4) <= DUpdateWireIns; wait for 1 ps;
      hi_in(1) <= '1'; wait for 1 ps;
      wait until (rising_edge(hi_clk)); hi_in(7 downto 4) <= DNOP; wait for 1 ps;
      for i in 0 to 31 loop
        hi_dataout <= WireIns(i); wait for 1 ps; wait until (rising_edge(hi_clk)); wait for 1 ps;
      end loop;
      wait until (hi_out(0) = '0'); wait for 1 ps; 
    end procedure UpdateWireIns;
     
    -----------------------------------------------------------------------
    -- UpdateWireOuts
    -----------------------------------------------------------------------
    procedure UpdateWireOuts is
      variable i : integer := 0;
    begin
      wait until (rising_edge(hi_clk)); hi_in(7 downto 4) <= DUpdateWireOuts; wait for 1 ps;
      wait until (rising_edge(hi_clk)); hi_in(7 downto 4) <= DNOP; wait for 1 ps;
      wait until (rising_edge(hi_clk)); hi_in(1) <= '0'; wait for 1 ps;
      wait until (rising_edge(hi_clk)); wait until (rising_edge(hi_clk)); wait for 1 ps;
      for i in 0 to 31 loop
        wait until (rising_edge(hi_clk)); WireOuts(i) := hi_inout; wait for 1 ps;
      end loop;
      wait until (hi_out(0) = '0'); wait for 1 ps;
    end procedure UpdateWireOuts;
  
    -----------------------------------------------------------------------
    -- ActivateTriggerIn
    -----------------------------------------------------------------------
    procedure ActivateTriggerIn (
      ep  : in  std_logic_vector(7 downto 0);
      bit : in  integer) is 
      
      variable tmp_slv4 :     std_logic_vector(3 downto 0);
    begin
      tmp_slv4 := CONV_std_logic_vector(bit, 4);
      wait until (rising_edge(hi_clk)); hi_in(7 downto 4) <= DActivateTriggerIn;
      hi_in(1) <= '1';
      hi_dataout <= (x"00" & ep);
      wait until (rising_edge(hi_clk)); hi_in(7 downto 4) <= DNOP;
      hi_dataout <= SHL(x"0001", tmp_slv4);
      wait until (rising_edge(hi_clk)); hi_dataout <= x"0000";
      wait until (hi_out(0) = '0');
    end procedure ActivateTriggerIn;
  
    -----------------------------------------------------------------------
    -- UpdateTriggerOuts
    -----------------------------------------------------------------------
    procedure UpdateTriggerOuts is
      variable i: integer := 0;
    begin
      wait until (rising_edge(hi_clk)); hi_in(7 downto 4) <= DUpdateTriggerOuts;
      wait until (rising_edge(hi_clk)); hi_in(7 downto 4) <= DNOP;
      wait until (rising_edge(hi_clk)); hi_in(1) <= '0';
      wait until (rising_edge(hi_clk)); wait until (rising_edge(hi_clk));
      wait until (rising_edge(hi_clk));
      
      for i in 0 to (UPDATE_TO_READOUT_CLOCKS-1) loop
          wait until (rising_edge(hi_clk));  
      end loop;
      
      for i in 0 to 31 loop
        wait until (rising_edge(hi_clk)); Triggered(i) := hi_inout;
      end loop;
      wait until (hi_out(0) = '0');
    end procedure UpdateTriggerOuts;
  
    -----------------------------------------------------------------------
    -- WriteToPipeIn
    -----------------------------------------------------------------------
    procedure WriteToPipeIn (
      ep      : in  std_logic_vector(7 downto 0);
      length  : in  integer) is
  
      variable len, i, j, k, blockSize : integer;
      variable tmp_slv8                : std_logic_vector(7 downto 0);
      variable tmp_slv32               : std_logic_vector(31 downto 0);
    begin
      len := (length / 2); j := 0; k := 0; blockSize := 1024;
      tmp_slv8 := CONV_std_logic_vector(BlockDelayStates, 8);
      tmp_slv32 := CONV_std_logic_vector(len, 32);
      wait until (rising_edge(hi_clk)); hi_in(1) <= '1';
      hi_in(7 downto 4) <= DWriteToPipeIn;
      hi_dataout <= (tmp_slv8 & ep);
      wait until (rising_edge(hi_clk)); hi_in(7 downto 4) <= DNOP;
      hi_dataout <= tmp_slv32(15 downto 0);
      wait until (rising_edge(hi_clk));
      hi_dataout <= tmp_slv32(31 downto 16);
      for i in 0 to len - 1 loop
        wait until (rising_edge(hi_clk));
        hi_dataout(7 downto 0) <= pipeIn(i*2);
        hi_dataout(15 downto 8) <= pipeIn((i*2)+1);
        j := j + 2;
        if (j = blockSize) then
          for k in 0 to BlockDelayStates - 1 loop
            wait until (rising_edge(hi_clk));
          end loop;
          j := 0;
        end if;
      end loop;
      wait until (hi_out(0) = '0');
    end procedure WriteToPipeIn;
  
    -----------------------------------------------------------------------
    -- ReadFromPipeOut
    -----------------------------------------------------------------------
    procedure ReadFromPipeOut (
      ep     : in  std_logic_vector(7 downto 0);
      length : in  integer) is
      
      variable len, i, j, k, blockSize : integer;
      variable tmp_slv8                : std_logic_vector(7 downto 0);
      variable tmp_slv32               : std_logic_vector(31 downto 0);
    begin
      len := (length / 2); j := 0; blockSize := 1024;
      tmp_slv8 := CONV_std_logic_vector(BlockDelayStates, 8);
      tmp_slv32 := CONV_std_logic_vector(len, 32);
      wait until (rising_edge(hi_clk)); hi_in(1) <= '1';
      hi_in(7 downto 4) <= DReadFromPipeOut;
      hi_dataout <= (tmp_slv8 & ep);
      wait until (rising_edge(hi_clk)); hi_in(7 downto 4) <= DNOP;
      hi_dataout <= tmp_slv32(15 downto 0);
      wait until (rising_edge(hi_clk));
      hi_dataout <= tmp_slv32(31 downto 16);
      wait until (rising_edge(hi_clk));
      hi_in(1) <= '0';
      for i in 0 to len - 1 loop
        wait until (rising_edge(hi_clk));
        pipeOut(i*2) := hi_inout(7 downto 0);
        pipeOut((i*2)+1) := hi_inout(15 downto 8);
        j := j + 2;
        if (j = blockSize) then
          for k in 0 to BlockDelayStates - 1 loop
            wait until (rising_edge(hi_clk));
          end loop;
          j := 0;
        end if;
      end loop;
      wait until (hi_out(0) = '0');
    end procedure ReadFromPipeOut;
  
    -----------------------------------------------------------------------
    -- WriteToBlockPipeIn
    -----------------------------------------------------------------------
    procedure WriteToBlockPipeIn (
      ep          : in std_logic_vector(7 downto 0);
      blockLength : in integer;
      length      : in integer) is
      
      variable len, i, j, k, blockSize, blockNum : integer;
      variable tmp_slv8                          : std_logic_vector(7 downto 0);
      variable tmp_slv16                         : std_logic_vector(15 downto 0);
      variable tmp_slv32                         : std_logic_vector(31 downto 0);
    begin
  
      len := (length/2); blockSize := (blockLength/2); j := 0; k := 0;
      blockNum := (len/blockSize);
      tmp_slv8 := CONV_std_logic_vector(BlockDelayStates, 8);
      tmp_slv32 := CONV_std_logic_vector(len, 32);
      wait until (rising_edge(hi_clk)); hi_in(1) <= '1';
      hi_in(7 downto 4) <= DWriteToBlockPipeIn;
      hi_dataout <= (tmp_slv8 & ep);
      wait until (rising_edge(hi_clk)); hi_in(7 downto 4) <= DNOP;
      hi_dataout <= tmp_slv32(15 downto 0);
      wait until (rising_edge(hi_clk)); hi_dataout <= tmp_slv32(31 downto 16);
      tmp_slv16 := CONV_std_logic_vector(blockSize, 16);
      wait until (rising_edge(hi_clk)); hi_dataout <= tmp_slv16;
      wait until (rising_edge(hi_clk));
      tmp_slv16 := (CONV_std_logic_vector(PostReadyDelay, 8) & CONV_std_logic_vector(ReadyCheckDelay, 8));
      hi_dataout <= tmp_slv16;
      for i in 1 to blockNum loop
        while (hi_out(0) = '1') loop wait until (rising_edge(hi_clk)); end loop;
        while (hi_out(0) = '0') loop wait until (rising_edge(hi_clk)); end loop;
        wait until (rising_edge(hi_clk)); wait until (rising_edge(hi_clk));
        for j in 1 to blockSize loop
          hi_dataout(7 downto 0) <= pipeIn(k);
          hi_dataout(15 downto 8) <= pipeIn(k+1);
          wait until (rising_edge(hi_clk)); k:=k+2;
        end loop;
        for j in 1 to BlockDelayStates loop 
          wait until (rising_edge(hi_clk)); 
        end loop;
      end loop;
      wait until (hi_out(0) = '0');
    end procedure WriteToBlockPipeIn;
  
    -----------------------------------------------------------------------
    -- ReadFromBlockPipeOut
    -----------------------------------------------------------------------
    procedure ReadFromBlockPipeOut (
      ep          : in std_logic_vector(7 downto 0);
      blockLength : in integer;
      length      : in integer) is
      
      variable len, i, j, k, blockSize, blockNum : integer;
      variable tmp_slv8                          : std_logic_vector(7 downto 0);
      variable tmp_slv16                         : std_logic_vector(15 downto 0);
      variable tmp_slv32                         : std_logic_vector(31 downto 0);
    begin
      len := (length/2); blockSize := (blockLength/2); j := 0; k := 0;
      blockNum := (len/blockSize);
      tmp_slv8 := CONV_std_logic_vector(BlockDelayStates, 8);
      tmp_slv32 := CONV_std_logic_vector(len, 32);
      wait until (rising_edge(hi_clk));
      hi_in(1) <= '1';
      hi_in(7 downto 4) <= DReadFromBlockPipeOut;
      hi_dataout <= (tmp_slv8 & ep);
      wait until (rising_edge(hi_clk)); hi_in(7 downto 4) <= DNOP;
      hi_dataout <= tmp_slv32(15 downto 0);
      wait until (rising_edge(hi_clk)); hi_dataout <= tmp_slv32(31 downto 16);
      tmp_slv16 := CONV_std_logic_vector(blockSize, 16);
      wait until (rising_edge(hi_clk)); hi_dataout <= tmp_slv16;
      wait until (rising_edge(hi_clk));
      tmp_slv16 := (CONV_std_logic_vector(PostReadyDelay, 8) & CONV_std_logic_vector(ReadyCheckDelay, 8));
      hi_dataout <= tmp_slv16;
      wait until (rising_edge(hi_clk)); hi_in(1) <= '0';
      for i in 1 to blockNum loop
        while (hi_out(0) = '1') loop wait until (rising_edge(hi_clk)); end loop;
        while (hi_out(0) = '0') loop wait until (rising_edge(hi_clk)); end loop;
        wait until (rising_edge(hi_clk)); wait until (rising_edge(hi_clk));
        for j in 1 to blockSize loop
          pipeOut(k) := hi_inout(7 downto 0); pipeOut(k+1) := hi_inout(15 downto 8);
          wait until (rising_edge(hi_clk)); k:=k+2;
        end loop;
        for j in 1 to BlockDelayStates loop wait until (rising_edge(hi_clk)); end loop;
      end loop;
      wait until (hi_out(0) = '0');
    end procedure ReadFromBlockPipeOut;




-- wireInLines unpacked:
-- [    | reloadCoef | runFIRFilter | run_mac | load_ram | rst ]
-- [    |    4       |    3         |      2  |   1      |  0  ]

   -- Stimulus process
   
   begin    


    FrontPanelReset;

      
      -- hold reset state for 100 ns.
      wait for 100 ns;  

      wait for clk1_period*10;
      report "Starting Simulation...";

      decimFactor <= 4;

      report "Pump the reset line...";
      -- set rst high:
      wireInLines <= x"0001"; wait until (rising_edge(clk1));
      SetWireInValue(x"00",wireInLines,x"ffff");
      UpdateWireIns;


      wireInLines <= x"0000"; wait until (rising_edge(clk1));
      SetWireInValue(x"00",wireInLines,x"ffff");
      UpdateWireIns;

      wait for clk1_period*10;

      -- load_ram high:
      wireInLines <= x"0002"; wait until (rising_edge(clk1));
      SetWireInValue(x"00",wireInLines,x"ffff");
      UpdateWireIns;
      report "Writing coefficients to block ram...";
      for i in 0 to windowSize loop
        windowCoef <= myCoef(i); wait until (rising_edge(clk1)); 
        SetWireInValue(x"07",std_logic_vector(conv_unsigned(i,16)),x"ffff");
        SetWireInValue(x"05",windowCoef(31 downto 16),x"ffff");
        SetWireInValue(x"06",windowCoef(15 downto 0),x"ffff");
        UpdateWireIns;
        ActivateTriggerIn(x"40",0);
        report "Address: " & integer'image(i);
      end loop;

      report "Writing inputSignal to wireIn...";
      for i in 0 to inputSize loop
        inputSignal <= myCosine(i); wait until (rising_edge(clk1)); 
        SetWireInValue(x"03",std_logic_vector(conv_unsigned(i,16)),x"ffff");
        SetWireInValue(x"02",inputSignal,x"ffff");
        UpdateWireIns;
        ActivateTriggerIn(x"40",0);
        report "Address: " & integer'image(i);
      end loop;

  
      wireInLines <= x"0000"; wait until (rising_edge(clk1));
      SetWireInValue(x"00",wireInLines,x"ffff");
      UpdateWireIns;

      -- runFilter high:
      wireInLines <= x"000C"; wait until (rising_edge(clk1));
      SetWireInValue(x"00",wireInLines,x"ffff");
      UpdateWireIns;
      report "Set Phase Increment for NCO...";
      phaseInc <= x"147A"; wait until (rising_edge(clk1));
      SetWireInValue(x"01",phaseInc,x"ffff");
      UpdateWireIns;      

      -- wait for 13 us;

      slow_clk <= (others => '0'); 

      report "Read data back from wireouts...";
      for i in 0 to windowSize loop
        -- slow_clk <= not slow_clk;
        -- SetWireInValue(x"08",slow_clk,x"ffff");
        SetWireInValue(x"04",std_logic_vector(conv_unsigned(i,16)),x"ffff"); wait for 1 ps;
        UpdateWireIns;
        report "Address: " & integer'image(i);
        UpdateWireOuts;
        acc_padRe2(63 downto 48) <= GetWireOutValue(x"20"); wait until (rising_edge(hi_clk)); -- wait for 1 ps; 
        acc_padRe2(47 downto 32) <= GetWireOutValue(x"21");  wait until (rising_edge(hi_clk)); -- wait for 1 ps; 
        acc_padRe2(31 downto 16) <= GetWireOutValue(x"22");  wait until (rising_edge(hi_clk)); -- wait for 1 ps; 
        acc_padRe2(15 downto 0) <= GetWireOutValue(x"23");  wait until (rising_edge(hi_clk)); -- wait for 1 ps; 

        acc_padIm2(63 downto 48) <= GetWireOutValue(x"24");  wait until (rising_edge(hi_clk)); -- wait for 1 ps; 
        acc_padIm2(47 downto 32) <= GetWireOutValue(x"25");  wait until (rising_edge(hi_clk)); -- wait for 1 ps; 
        acc_padIm2(31 downto 16) <= GetWireOutValue(x"26");  wait until (rising_edge(hi_clk)); -- wait for 1 ps; 
        acc_padIm2(15 downto 0) <= GetWireOutValue(x"27");  wait until (rising_edge(hi_clk)); -- wait for 1 ps; 
        acc <= acc_padIm2(49 downto 0) & acc_padRe2(49 downto 0); wait until (rising_edge(hi_clk));

      end loop;

      wireInLines <= x"0000"; wait until (rising_edge(clk1));
      SetWireInValue(x"00",wireInLines,x"ffff");
      UpdateWireIns;
      

      report "Finished Processing.";


     wait;
   end process;

end behavior;
